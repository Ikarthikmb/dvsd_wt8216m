// 8 bit Multiplier
// 
// A           0000 0000
// B           0000 0000
// -----------------------
//             0000 0000
//           0 0000 000
//          00 0000 00
//         000 0000 0
//        0000 0000
//      0 0000 000
//     00 0000 00
//    000 0000 0
// -----------------------
// M 0000 0000 0000 0000
// -----------------------

module dvsd_8216m9(
	input  [7:0] A,
	input  [7:0] B,
	output [15:0] M
	);
	
	assign M = A * B;
endmodule

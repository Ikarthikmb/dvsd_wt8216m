// ==============================================================
// 
// AND Gate
// 
// ==============================================================

module and1b(
  input a1,
  input a2,
  output y
);

  assign y = a1 & a2;
  
endmodule
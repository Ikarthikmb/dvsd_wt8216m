// 4:2 Compressor

// `include "cmos_inverter.v"

module compressor4to2(
	input a0,
	input a1,
	input a2,
	input a3,
	output sout,
	output cout
);
	supply0 GND;
	supply1 PWR;

	//SUM Logic
	
	//CARRY Logic
	
endmodule

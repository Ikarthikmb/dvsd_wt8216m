* SPICE3 file created from dvsd_8216m9.ext - technology: sky130A

.subckt dvsd_8216m9 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] B[0] B[1] B[2] B[3] B[4]
+ B[5] B[6] B[7] M[0] M[10] M[11] M[12] M[13] M[14] M[15] M[1] M[2] M[3] M[4] M[5]
+ M[6] M[7] M[8] M[9] VGND VPWR
C0 _567_/B _571_/a_250_297# 0.13fF
C1 _480_/Y _542_/A 0.16fF
C2 _375_/a_79_199# _375_/a_448_47# 0.13fF
C3 _566_/A _570_/B 0.03fF
C4 B[7] _574_/X 0.07fF
C5 _487_/a_78_199# _452_/X 0.13fF
C6 B[1] _584_/A 0.12fF
C7 _396_/X _392_/Y 0.11fF
C8 _542_/C _505_/a_80_21# 0.09fF
C9 _441_/a_78_199# _454_/X 0.12fF
C10 _548_/a_489_413# _546_/X 0.15fF
C11 _634_/a_27_413# _368_/A 0.09fF
C12 _508_/a_77_199# _508_/a_539_297# 0.06fF
C13 _316_/a_381_47# _316_/a_558_47# 0.32fF
C14 _322_/A VPWR 1.38fF
C15 _557_/B _558_/a_323_297# 0.13fF
C16 _626_/a_109_47# _626_/Y 0.50fF
C17 _543_/A _515_/A 0.21fF
C18 _358_/a_109_47# _485_/A 0.04fF
C19 _542_/C _443_/B 1.04fF
C20 _613_/X _589_/a_489_413# 0.13fF
C21 _611_/a_109_297# _611_/X 0.03fF
C22 _616_/A _530_/X 0.28fF
C23 _630_/X _363_/B 0.01fF
C24 B[0] _514_/B 0.28fF
C25 _583_/X _580_/B 0.50fF
C26 _516_/A _542_/A 0.03fF
C27 _539_/A _542_/A 0.85fF
C28 _569_/A _612_/Y 0.03fF
C29 _593_/A _598_/A 0.11fF
C30 _440_/X _460_/a_489_413# 0.07fF
C31 _587_/A A[6] 0.08fF
C32 _614_/a_489_413# VPWR 0.39fF
C33 _574_/X _574_/a_81_21# 0.24fF
C34 _340_/A _381_/B 0.16fF
C35 _469_/A _521_/X 0.94fF
C36 _352_/a_222_93# _314_/X 0.03fF
C37 _539_/a_150_297# _442_/A 0.01fF
C38 _556_/Y _582_/a_27_47# 0.01fF
C39 _627_/A _586_/a_505_21# 0.21fF
C40 _455_/X _389_/a_27_47# 0.10fF
C41 _458_/X _437_/X 0.15fF
C42 _557_/Y VPWR 2.31fF
C43 VPWR _483_/a_250_297# 0.74fF
C44 _602_/A VPWR 1.99fF
C45 B[7] _549_/a_76_199# 0.06fF
C46 _337_/a_150_297# _338_/X 0.02fF
C47 _457_/X VPWR 1.15fF
C48 _545_/Y _546_/a_489_413# 0.14fF
C49 _588_/A _381_/B 0.08fF
C50 _610_/A _621_/a_292_297# 0.02fF
C51 _433_/Y _540_/a_93_21# 0.05fF
C52 _419_/a_226_47# _419_/X 0.05fF
C53 _443_/A _441_/a_215_47# 0.01fF
C54 _448_/B _542_/D 1.35fF
C55 _551_/X _530_/X 1.43fF
C56 _413_/X _419_/a_226_47# 0.24fF
C57 _556_/Y _558_/a_323_297# 0.02fF
C58 _557_/A _558_/a_227_47# 0.02fF
C59 _467_/Y VPWR 3.46fF
C60 _620_/a_489_413# _619_/Y 0.14fF
C61 _627_/X _608_/X 0.09fF
C62 _433_/Y _621_/X 0.75fF
C63 _498_/Y _527_/Y 0.31fF
C64 _461_/a_493_297# VPWR 0.01fF
C65 _566_/A _381_/B 1.58fF
C66 _510_/A _387_/a_215_47# 0.16fF
C67 _491_/a_76_199# _491_/X 0.22fF
C68 _612_/Y _627_/D 0.35fF
C69 _627_/C _627_/a_27_297# 0.45fF
C70 _329_/a_76_199# _352_/a_448_47# 0.00fF
C71 _580_/B _580_/a_68_297# 0.43fF
C72 _446_/X _469_/X 0.03fF
C73 _544_/A _561_/A 1.41fF
C74 _586_/S _621_/X 0.00fF
C75 _458_/X _439_/a_76_199# 0.07fF
C76 _416_/a_215_47# _418_/A 0.15fF
C77 _417_/A _417_/a_27_47# 0.43fF
C78 _504_/a_77_199# _390_/B 0.01fF
C79 _453_/X _453_/a_93_21# 0.13fF
C80 _519_/A _519_/C 0.28fF
C81 _417_/D _480_/A 0.13fF
C82 _336_/a_215_47# _328_/A 0.11fF
C83 _495_/a_226_47# _497_/A 0.05fF
C84 _627_/X _627_/C 0.06fF
C85 input11/a_27_47# _485_/D 0.24fF
C86 B[7] _590_/a_150_297# 0.02fF
C87 _510_/A _393_/A 0.90fF
C88 _338_/a_544_297# _332_/X 0.04fF
C89 _595_/a_323_297# _566_/Y 0.03fF
C90 _540_/X _540_/a_93_21# 0.13fF
C91 _342_/X _352_/a_222_93# 0.13fF
C92 _412_/a_76_199# _408_/X 0.36fF
C93 _425_/a_76_199# _426_/B 0.22fF
C94 _500_/a_78_199# _497_/a_68_297# 0.00fF
C95 _547_/a_79_199# _547_/X 0.29fF
C96 _410_/B _485_/A 0.36fF
C97 _459_/X VPWR 0.76fF
C98 _563_/A _518_/X 0.03fF
C99 _581_/a_27_93# _581_/B 0.47fF
C100 _469_/a_62_47# _588_/A 0.14fF
C101 _361_/X _374_/X 0.34fF
C102 _432_/A _371_/A 0.35fF
C103 _577_/a_556_47# _390_/D 0.02fF
C104 _351_/A _351_/X 0.07fF
C105 _574_/X VPWR 3.69fF
C106 _503_/A VPWR 5.69fF
C107 _543_/A _469_/a_664_47# 0.01fF
C108 _467_/Y _501_/Y 1.34fF
C109 _417_/D _481_/A 0.02fF
C110 _428_/a_384_47# _427_/Y 0.01fF
C111 _578_/a_78_199# VPWR 0.61fF
C112 _623_/a_226_47# _433_/Y 0.11fF
C113 _386_/a_664_47# _515_/A 0.07fF
C114 _631_/Y _316_/a_381_47# 0.08fF
C115 _626_/Y _559_/X 0.03fF
C116 output21/a_27_47# _626_/a_109_47# 0.01fF
C117 _544_/a_664_47# _503_/A 0.01fF
C118 _615_/a_493_297# _593_/Y 0.08fF
C119 _417_/D _633_/Y 0.05fF
C120 _387_/a_493_297# _475_/A 0.02fF
C121 _347_/A _481_/A 0.05fF
C122 _548_/a_76_199# _548_/a_489_413# 0.12fF
C123 _613_/a_77_199# _590_/A 0.03fF
C124 _419_/a_76_199# _452_/A 0.10fF
C125 _359_/a_68_297# _383_/X 0.14fF
C126 _391_/A _420_/X 0.04fF
C127 _474_/A _473_/a_227_47# 0.04fF
C128 VPWR _606_/A 4.00fF
C129 M[0] _554_/A 0.09fF
C130 _599_/A _575_/X 0.01fF
C131 _416_/a_292_297# _561_/A 0.04fF
C132 _350_/a_109_297# _350_/C 0.08fF
C133 VPWR _609_/a_209_297# 0.45fF
C134 _357_/a_27_47# _509_/A 0.01fF
C135 _347_/A _633_/Y 0.08fF
C136 _337_/B _631_/B 0.40fF
C137 _634_/a_27_413# _370_/A 0.37fF
C138 _586_/S _586_/a_76_199# 0.65fF
C139 _340_/A _542_/A 0.12fF
C140 _603_/Y output17/a_27_47# 0.01fF
C141 VPWR _427_/A 2.16fF
C142 _504_/a_323_297# _471_/Y 0.05fF
C143 _433_/a_481_47# _432_/X 0.09fF
C144 output32/a_27_47# M[9] 0.44fF
C145 _498_/Y _531_/A 0.10fF
C146 _606_/Y _606_/A 1.10fF
C147 _468_/a_215_47# _436_/X 0.03fF
C148 _626_/Y _465_/X 0.03fF
C149 _485_/D _484_/a_78_199# 0.14fF
C150 _507_/Y _539_/X 0.23fF
C151 _588_/A _593_/A 0.36fF
C152 _590_/B _622_/C 0.26fF
C153 _610_/A _624_/a_489_47# 0.07fF
C154 _497_/A _494_/X 0.01fF
C155 _635_/a_27_413# _635_/a_300_297# 0.04fF
C156 _626_/Y _616_/B 0.85fF
C157 _331_/a_27_47# _351_/a_27_53# 0.01fF
C158 _474_/A _476_/a_250_297# 0.03fF
C159 _503_/A _559_/a_539_297# 0.08fF
C160 _456_/a_489_413# VPWR 0.39fF
C161 _549_/a_76_199# VPWR 0.50fF
C162 _390_/a_27_47# VPWR 0.80fF
C163 _453_/a_93_21# _542_/D 0.36fF
C164 _525_/a_226_47# _523_/X 0.29fF
C165 _424_/a_226_47# VPWR 0.16fF
C166 _359_/A _447_/B 0.15fF
C167 _566_/A _542_/A 0.35fF
C168 _587_/A _472_/Y 0.21fF
C169 _465_/X _467_/a_109_47# 0.20fF
C170 _568_/a_227_47# _433_/Y 0.07fF
C171 _444_/Y _390_/B 0.27fF
C172 _567_/B A[3] 0.05fF
C173 _351_/A _419_/X 0.11fF
C174 _563_/A _520_/X 0.28fF
C175 _542_/B _478_/a_27_47# 0.36fF
C176 _455_/X _631_/Y 0.30fF
C177 _423_/X _461_/X 0.02fF
C178 _591_/Y B[7] 0.11fF
C179 _516_/A _519_/X 0.12fF
C180 _382_/B _420_/X 0.06fF
C181 _559_/X _381_/B 0.03fF
C182 _602_/Y _554_/B 0.73fF
C183 _454_/a_76_199# _449_/A 0.02fF
C184 _631_/Y _509_/A 0.23fF
C185 _359_/A _376_/a_68_297# 0.03fF
C186 _471_/Y VPWR 2.30fF
C187 _326_/A _350_/C 0.48fF
C188 _330_/A _363_/A 0.03fF
C189 _627_/A _520_/X 0.37fF
C190 _427_/A _501_/Y 0.11fF
C191 _538_/Y _539_/X 0.55fF
C192 _544_/A VPWR 5.80fF
C193 _627_/A _590_/A 0.30fF
C194 _568_/a_227_297# _546_/X 0.03fF
C195 _355_/A _316_/a_381_47# 0.01fF
C196 _330_/A _420_/X 0.79fF
C197 _381_/C _520_/a_489_413# 0.09fF
C198 _485_/a_27_47# _485_/A 0.37fF
C199 _536_/Y _539_/A 0.01fF
C200 _510_/A _433_/Y 1.53fF
C201 _544_/A _544_/a_664_47# 0.07fF
C202 _381_/C _519_/A 0.15fF
C203 _474_/A _509_/Y 0.01fF
C204 B[2] _576_/X 0.53fF
C205 _390_/D _538_/A 0.50fF
C206 _487_/a_78_199# _447_/B 0.01fF
C207 _379_/a_78_199# _419_/a_76_199# 0.01fF
C208 _318_/a_27_47# _563_/A 0.04fF
C209 _440_/X _459_/a_556_47# 0.02fF
C210 _423_/X _407_/a_27_47# 0.00fF
C211 _589_/a_76_199# _590_/B 0.23fF
C212 _447_/B _367_/C 0.03fF
C213 _404_/a_558_47# _442_/D 0.10fF
C214 VPWR _446_/a_93_21# 0.36fF
C215 _584_/A _547_/X 0.03fF
C216 _542_/D _514_/B 0.27fF
C217 A[6] _484_/a_78_199# 0.05fF
C218 _504_/a_227_47# _436_/X 0.01fF
C219 _531_/B _558_/X 0.17fF
C220 _433_/Y _485_/D 0.02fF
C221 _571_/a_93_21# _381_/B 0.30fF
C222 _391_/B VPWR 1.38fF
C223 _452_/A _628_/Y 1.02fF
C224 _585_/B _593_/Y 0.05fF
C225 _444_/Y _471_/A 0.03fF
C226 VPWR _504_/X 4.33fF
C227 _467_/Y _531_/C 0.03fF
C228 _621_/a_78_199# _621_/a_292_297# 0.03fF
C229 _375_/a_79_199# _519_/A 0.17fF
C230 _466_/a_215_47# _466_/X 0.01fF
C231 _566_/Y VPWR 2.59fF
C232 _594_/a_109_297# _595_/X 0.09fF
C233 B[2] _618_/A 0.52fF
C234 _539_/X _486_/X 0.24fF
C235 _587_/A _437_/X 0.33fF
C236 _406_/A _458_/X 0.09fF
C237 _502_/a_215_47# _492_/X 0.11fF
C238 _567_/a_109_297# VPWR 0.01fF
C239 _545_/Y _610_/A 1.19fF
C240 _416_/a_292_297# VPWR 0.01fF
C241 _437_/X _439_/a_489_413# 0.26fF
C242 _455_/X _490_/a_78_199# 0.15fF
C243 _397_/a_76_199# _397_/a_226_47# 0.49fF
C244 _417_/D _515_/Y 0.07fF
C245 _436_/A _412_/a_76_199# 0.04fF
C246 _386_/A _470_/a_209_297# 0.07fF
C247 _485_/D _540_/X 0.04fF
C248 _433_/Y _483_/X 0.03fF
C249 _454_/X _519_/C 0.80fF
C250 _445_/A _387_/a_292_297# 0.08fF
C251 _447_/X _449_/A 0.73fF
C252 _487_/X _538_/Y 0.33fF
C253 _347_/A _515_/Y 0.16fF
C254 _382_/X _452_/A 1.47fF
C255 _343_/a_489_413# _329_/X 0.17fF
C256 _605_/a_209_297# _604_/a_209_297# 0.01fF
C257 _452_/A _452_/X 0.23fF
C258 _491_/X _524_/X 0.05fF
C259 _423_/a_78_199# _423_/a_292_297# 0.03fF
C260 _426_/A _432_/X 0.30fF
C261 _568_/a_77_199# _536_/Y 0.02fF
C262 _406_/B _390_/B 0.03fF
C263 _570_/B _530_/X 0.27fF
C264 _441_/a_78_199# VPWR 0.64fF
C265 _330_/A _374_/X 0.37fF
C266 _626_/Y _530_/X 0.03fF
C267 _587_/A _590_/B 0.47fF
C268 _587_/A _439_/a_76_199# 0.05fF
C269 _439_/a_76_199# _439_/a_489_413# 0.12fF
C270 _562_/a_78_199# _584_/A 0.42fF
C271 _493_/a_78_199# _493_/a_292_297# 0.03fF
C272 B[2] _549_/X 0.03fF
C273 _386_/A _547_/X 0.30fF
C274 _503_/a_62_47# _503_/a_381_47# 0.08fF
C275 _629_/B _371_/B 0.22fF
C276 _338_/a_79_199# _338_/X 0.29fF
C277 _540_/X _483_/X 0.05fF
C278 _614_/a_556_47# _612_/Y 0.02fF
C279 _563_/B _449_/A 0.20fF
C280 _439_/X _458_/X 0.36fF
C281 _508_/a_77_199# _507_/Y 0.44fF
C282 _591_/Y VPWR 3.33fF
C283 _590_/B _612_/A 0.31fF
C284 _420_/X _421_/a_76_199# 0.26fF
C285 _613_/a_77_199# _503_/A 0.00fF
C286 _596_/a_489_413# _600_/a_27_297# 0.01fF
C287 _350_/a_277_297# _442_/B 0.01fF
C288 _429_/a_76_199# B[5] 0.02fF
C289 _632_/a_215_47# _475_/A 0.12fF
C290 _534_/a_80_21# _381_/B 0.26fF
C291 _543_/B _542_/C 0.08fF
C292 _537_/a_227_297# _535_/Y 0.01fF
C293 _627_/D _621_/a_292_297# 0.02fF
C294 _587_/a_27_47# VPWR 0.50fF
C295 A[6] _433_/Y 0.05fF
C296 _419_/X _519_/A 0.54fF
C297 _380_/A _326_/A 0.03fF
C298 _621_/a_215_47# _591_/A 0.11fF
C299 _629_/A _363_/B 0.05fF
C300 _376_/X _383_/X 0.84fF
C301 _633_/Y _595_/X 0.03fF
C302 _328_/A _475_/A 0.25fF
C303 _616_/B _593_/A 0.66fF
C304 _487_/X _486_/X 4.08fF
C305 _378_/A _485_/D 0.09fF
C306 _625_/Y _590_/B 0.18fF
C307 _420_/X _442_/B 0.20fF
C308 _587_/A _506_/Y 0.21fF
C309 _539_/a_68_297# _539_/a_150_297# 0.02fF
C310 _538_/Y _570_/A 0.53fF
C311 _605_/a_80_21# VPWR 0.36fF
C312 _417_/D _585_/B 0.42fF
C313 _513_/A _487_/X 0.03fF
C314 input3/a_841_47# _616_/Y 0.02fF
C315 input3/a_664_47# _616_/A 0.00fF
C316 _462_/a_76_199# _462_/a_489_413# 0.12fF
C317 _569_/Y _621_/X 0.09fF
C318 _573_/A VPWR 2.20fF
C319 _408_/B _408_/X 0.01fF
C320 _623_/a_489_413# _628_/Y 0.03fF
C321 _474_/Y VPWR 0.99fF
C322 B[0] _562_/a_215_47# 0.02fF
C323 _524_/a_78_199# _524_/a_215_47# 0.26fF
C324 output24/a_27_47# _627_/D 0.00fF
C325 B[0] _472_/B 0.38fF
C326 _480_/Y _539_/A 0.11fF
C327 _630_/X _398_/a_76_199# 0.07fF
C328 _544_/a_62_47# _544_/a_558_47# 0.03fF
C329 _530_/X _381_/B 1.91fF
C330 _442_/B _411_/A 0.08fF
C331 _619_/a_27_47# VPWR 0.04fF
C332 _375_/a_222_93# _447_/B 0.00fF
C333 _542_/B _411_/A 0.09fF
C334 _327_/a_78_199# _367_/C 0.30fF
C335 _378_/a_62_47# _542_/D 0.12fF
C336 _513_/A _381_/C 2.27fF
C337 _540_/a_93_21# _540_/a_346_47# 0.05fF
C338 _627_/A _503_/A 2.59fF
C339 _445_/A _350_/C 1.49fF
C340 _523_/X _492_/a_489_413# 0.01fF
C341 _527_/A _530_/X 0.18fF
C342 _619_/a_27_47# _606_/Y 0.08fF
C343 _516_/A _539_/A 0.29fF
C344 _579_/X M[0] 0.05fF
C345 _417_/A _369_/a_556_47# 0.05fF
C346 _480_/A _410_/C 0.17fF
C347 _444_/A VPWR 3.09fF
C348 _375_/a_222_93# _376_/a_68_297# 0.01fF
C349 _411_/a_150_297# _510_/A 0.01fF
C350 _328_/X _442_/B 0.59fF
C351 VPWR B[5] 4.49fF
C352 _404_/a_62_47# _503_/A 0.31fF
C353 _592_/a_113_297# _593_/A 0.22fF
C354 _635_/Y output26/a_27_47# 0.40fF
C355 _549_/X _551_/a_226_47# 0.26fF
C356 _550_/X _551_/a_489_413# 0.14fF
C357 _570_/A _486_/X 0.68fF
C358 _390_/D _390_/B 1.99fF
C359 _417_/D _447_/X 0.05fF
C360 _381_/C _454_/X 0.99fF
C361 _612_/Y _601_/A 0.10fF
C362 _350_/C _350_/B 0.28fF
C363 _464_/A _466_/X 1.51fF
C364 _574_/X _548_/X 0.17fF
C365 _536_/a_109_297# _585_/B 0.02fF
C366 _386_/a_558_47# _570_/A 0.08fF
C367 _381_/C _334_/a_27_47# 0.37fF
C368 _575_/X _547_/X 0.01fF
C369 _335_/a_381_47# _335_/a_558_47# 0.32fF
C370 _542_/C _486_/X 0.04fF
C371 _418_/X _367_/C 0.14fF
C372 _445_/A _367_/C 0.39fF
C373 _378_/A A[6] 0.03fF
C374 _336_/a_493_297# _519_/A 0.05fF
C375 _557_/A _604_/X 0.05fF
C376 _404_/a_381_47# _609_/a_80_21# 0.03fF
C377 _534_/a_80_21# _542_/A 0.00fF
C378 _447_/a_68_297# output32/a_27_47# 0.00fF
C379 _542_/C _386_/a_558_47# 0.10fF
C380 _481_/A _410_/C 0.73fF
C381 _361_/a_556_47# _361_/X 0.02fF
C382 _513_/A _542_/C 0.69fF
C383 _442_/B _374_/X 0.17fF
C384 _476_/a_584_47# _469_/X 0.02fF
C385 _343_/a_226_47# _369_/a_226_47# 0.02fF
C386 _615_/a_215_47# _594_/X 0.03fF
C387 _340_/A _340_/a_27_47# 0.37fF
C388 VPWR _394_/a_558_47# 0.24fF
C389 _368_/B _337_/X 0.21fF
C390 _410_/B _470_/a_209_297# 0.09fF
C391 _511_/a_250_297# _509_/A 0.03fF
C392 _469_/A _571_/a_250_297# 0.02fF
C393 _476_/X _490_/X 0.20fF
C394 _465_/a_27_297# VPWR 0.65fF
C395 _627_/C _449_/A 0.28fF
C396 _561_/A _519_/C 0.20fF
C397 _400_/a_209_297# _391_/B 0.03fF
C398 _519_/a_29_53# _563_/B 0.46fF
C399 input2/a_27_47# _390_/B 0.43fF
C400 _583_/X A[3] 0.03fF
C401 _417_/D _563_/B 0.39fF
C402 _537_/a_77_199# _539_/X 0.01fF
C403 _402_/a_27_47# _439_/a_489_413# 0.02fF
C404 _455_/X _447_/B 0.71fF
C405 _563_/D _420_/X 0.14fF
C406 _630_/a_226_47# _426_/A 0.16fF
C407 B[7] _519_/C 0.02fF
C408 A[6] _505_/a_80_21# 0.10fF
C409 _454_/X _316_/a_62_47# 0.14fF
C410 _559_/a_77_199# _559_/a_323_297# 0.05fF
C411 _411_/a_68_297# _475_/A 0.07fF
C412 _408_/a_68_297# _631_/B 0.08fF
C413 _381_/a_27_47# _485_/A 0.61fF
C414 _542_/C _454_/X 0.29fF
C415 _442_/B _329_/X 0.12fF
C416 _584_/a_68_297# _621_/X 0.08fF
C417 _546_/a_226_47# VPWR 0.07fF
C418 _544_/A _563_/A 0.03fF
C419 _568_/a_77_199# _435_/a_27_47# 0.02fF
C420 _494_/a_76_199# _495_/a_226_47# 0.01fF
C421 _626_/Y _467_/a_109_297# 0.04fF
C422 _387_/a_78_199# VPWR 0.61fF
C423 _472_/Y _433_/Y 0.03fF
C424 _375_/X _352_/X 0.10fF
C425 _583_/X M[15] 0.00fF
C426 _610_/A _624_/X 0.12fF
C427 _510_/X _631_/Y 0.25fF
C428 _549_/a_76_199# _548_/X 0.22fF
C429 _549_/a_226_47# _540_/X 0.25fF
C430 _511_/a_93_21# _631_/Y 0.04fF
C431 _577_/a_76_199# _580_/A 0.22fF
C432 _546_/a_226_47# _544_/a_664_47# 0.01fF
C433 _627_/A _471_/Y 1.11fF
C434 _527_/A _557_/B 0.03fF
C435 _440_/a_76_199# VPWR 0.46fF
C436 _530_/X _542_/A 0.15fF
C437 _596_/a_76_199# _599_/Y 0.00fF
C438 _423_/a_215_47# _383_/X 0.10fF
C439 _563_/D _411_/A 0.03fF
C440 A[2] _618_/Y 0.02fF
C441 _379_/a_78_199# _379_/a_292_297# 0.03fF
C442 _564_/A _621_/X 0.00fF
C443 _626_/Y _462_/X 0.17fF
C444 _385_/a_841_47# VPWR 0.41fF
C445 _515_/Y _518_/a_93_21# 0.30fF
C446 _469_/A _535_/Y 0.01fF
C447 _426_/B _464_/Y 0.01fF
C448 _516_/a_27_47# _520_/X 0.07fF
C449 _569_/A _545_/Y 0.09fF
C450 _465_/a_27_297# _501_/Y 0.01fF
C451 _380_/A _486_/B 0.13fF
C452 _584_/A _481_/A 1.03fF
C453 _342_/X B[5] 0.30fF
C454 _446_/a_93_21# _470_/a_80_21# 0.07fF
C455 _633_/Y _584_/A 0.03fF
C456 _520_/a_226_297# _518_/X 0.02fF
C457 _520_/a_76_199# _520_/a_226_47# 0.49fF
C458 _383_/a_76_199# _383_/a_226_47# 0.49fF
C459 _373_/Y _430_/X 0.16fF
C460 _428_/a_299_297# _426_/B 0.07fF
C461 _443_/A _443_/B 0.16fF
C462 _516_/A _479_/A 0.79fF
C463 _328_/B _328_/A 0.56fF
C464 _610_/A _622_/C 0.77fF
C465 _340_/A _539_/A 0.10fF
C466 _487_/X _537_/a_77_199# 0.12fF
C467 _479_/A _539_/A 0.24fF
C468 _516_/A _340_/A 1.51fF
C469 _406_/Y _462_/X 2.10fF
C470 _445_/A _380_/A 0.03fF
C471 _378_/A _418_/B 1.33fF
C472 _452_/A _447_/B 0.13fF
C473 _589_/a_489_413# A[3] 0.09fF
C474 _627_/A _504_/X 0.04fF
C475 VPWR _482_/X 0.75fF
C476 _475_/A _631_/Y 0.03fF
C477 _557_/A _531_/B 0.50fF
C478 _435_/a_27_47# _588_/A 0.10fF
C479 input16/a_27_47# _540_/X 0.00fF
C480 _439_/X _587_/A 0.30fF
C481 _526_/a_226_47# _527_/B 0.05fF
C482 _559_/a_227_47# _535_/Y 0.13fF
C483 _576_/a_556_47# _485_/D 0.02fF
C484 _355_/a_161_47# _563_/D 0.14fF
C485 _627_/A _566_/Y 2.03fF
C486 VPWR _430_/X 1.79fF
C487 _381_/B _514_/B 0.51fF
C488 _351_/A _631_/A 0.03fF
C489 _386_/A _480_/A 0.00fF
C490 _436_/A _408_/B 1.27fF
C491 VPWR _531_/a_109_297# 0.01fF
C492 _380_/A _350_/B 2.10fF
C493 _487_/X _561_/A 0.17fF
C494 _381_/C _627_/B 0.01fF
C495 _347_/A _322_/a_27_47# 0.02fF
C496 _494_/a_226_47# _468_/X 0.01fF
C497 _538_/Y _540_/a_93_21# 0.22fF
C498 _494_/a_76_199# _494_/X 0.34fF
C499 _363_/A _397_/X 0.12fF
C500 _452_/A _376_/a_68_297# 0.00fF
C501 _396_/a_250_297# _386_/X 0.13fF
C502 _385_/a_62_47# _385_/a_381_47# 0.08fF
C503 input12/a_381_47# input12/a_558_47# 0.32fF
C504 _585_/B _595_/X 0.01fF
C505 _381_/C _448_/a_150_297# 0.02fF
C506 _437_/X _433_/Y 0.56fF
C507 _579_/a_59_75# _579_/a_145_75# 0.02fF
C508 _335_/a_664_47# _510_/A 0.05fF
C509 _503_/a_381_47# _475_/A 0.01fF
C510 _474_/A _469_/X 0.23fF
C511 _633_/A _631_/B 0.07fF
C512 _479_/a_68_297# _479_/a_150_297# 0.02fF
C513 _371_/B output26/a_27_47# 0.02fF
C514 _541_/a_78_199# _541_/a_292_297# 0.03fF
C515 B[0] _517_/X 0.05fF
C516 _386_/A _481_/A 0.36fF
C517 _350_/B _384_/a_226_47# 0.11fF
C518 VPWR _519_/C 4.27fF
C519 _480_/A _483_/a_93_21# 0.02fF
C520 _381_/C _561_/A 0.16fF
C521 _417_/D _627_/C 0.08fF
C522 _386_/A _633_/Y 0.34fF
C523 _343_/a_226_297# VPWR 0.00fF
C524 _436_/A _436_/a_68_297# 0.32fF
C525 _448_/A _628_/Y 0.03fF
C526 _485_/a_27_47# _547_/X 0.01fF
C527 _331_/a_27_47# _363_/A 0.07fF
C528 _537_/a_77_199# _570_/A 0.24fF
C529 _381_/C B[7] 0.31fF
C530 _375_/X _436_/A 0.03fF
C531 _580_/A _579_/X 0.24fF
C532 _378_/a_664_47# VPWR 0.49fF
C533 _587_/A _442_/A 0.26fF
C534 _629_/B _433_/Y 0.01fF
C535 _408_/B _350_/X 0.10fF
C536 _419_/X _337_/A 0.03fF
C537 _540_/a_93_21# _486_/X 0.10fF
C538 _497_/A _527_/a_109_297# 0.04fF
C539 VPWR _539_/X 2.18fF
C540 B[1] _391_/A 0.21fF
C541 _483_/a_93_21# _481_/A 0.01fF
C542 _510_/A _519_/A 0.46fF
C543 _594_/a_27_297# _574_/X 0.02fF
C544 _416_/a_215_47# _324_/a_62_47# 0.05fF
C545 _463_/a_226_297# VPWR 0.00fF
C546 _350_/a_27_297# _350_/a_109_297# 0.02fF
C547 _530_/a_76_199# _530_/X 0.32fF
C548 _543_/a_109_297# _543_/B 0.04fF
C549 _513_/A _547_/a_544_297# 0.04fF
C550 _493_/X _468_/X 0.06fF
C551 _551_/X _554_/A 0.01fF
C552 _448_/A _452_/X 0.03fF
C553 _463_/a_76_199# _626_/Y 0.08fF
C554 _386_/X _480_/A 0.02fF
C555 _396_/X _386_/X 0.12fF
C556 _568_/a_539_297# _567_/B 0.02fF
C557 VPWR _556_/A 2.62fF
C558 _568_/a_77_199# _566_/A 0.31fF
C559 _469_/A A[3] 0.97fF
C560 _455_/X _418_/X 0.00fF
C561 _631_/Y _511_/X 2.76fF
C562 _442_/D _479_/B 0.01fF
C563 _416_/a_493_297# _378_/A 0.09fF
C564 _527_/Y _531_/B 0.02fF
C565 _506_/Y _433_/Y 0.03fF
C566 _623_/X _612_/Y 0.46fF
C567 _519_/A _485_/D 0.01fF
C568 _474_/Y _627_/A 0.14fF
C569 _537_/a_77_199# _535_/A 0.16fF
C570 _499_/a_81_21# VPWR 0.49fF
C571 _478_/A _472_/B 0.08fF
C572 _340_/A _479_/A 0.01fF
C573 _397_/X _374_/X 1.46fF
C574 _443_/B _446_/a_250_297# 0.02fF
C575 VPWR _432_/a_68_297# 0.26fF
C576 _427_/Y _426_/A 0.88fF
C577 _542_/A _514_/B 0.06fF
C578 _567_/B _520_/X 0.03fF
C579 _519_/X _530_/X 0.08fF
C580 _466_/a_215_47# _431_/X 0.03fF
C581 _466_/a_78_199# _428_/X 0.01fF
C582 _635_/Y _635_/a_27_413# 0.35fF
C583 VPWR _575_/a_215_47# 0.08fF
C584 _390_/B _631_/Y 0.17fF
C585 _411_/a_68_297# _471_/A 0.01fF
C586 _632_/a_292_297# VPWR 0.01fF
C587 _375_/X _350_/X 0.03fF
C588 _406_/A _393_/A 0.09fF
C589 _412_/a_226_47# _412_/X 0.05fF
C590 _587_/A _610_/A 0.52fF
C591 _585_/B _410_/C 0.65fF
C592 _386_/X _481_/A 0.17fF
C593 _559_/a_539_297# _539_/X 0.02fF
C594 _533_/a_323_297# _503_/A 0.07fF
C595 _463_/a_76_199# _406_/Y 0.34fF
C596 _610_/A _612_/A 1.25fF
C597 _610_/Y _590_/B 0.01fF
C598 _444_/A _470_/a_80_21# 0.00fF
C599 _386_/X _633_/Y 0.03fF
C600 _595_/X _572_/B 0.08fF
C601 _410_/a_27_47# _410_/a_109_47# 0.03fF
C602 _536_/Y _530_/X 0.10fF
C603 input5/a_62_47# input5/a_558_47# 0.03fF
C604 B[0] _442_/D 0.05fF
C605 _444_/Y _390_/D 0.13fF
C606 _327_/a_78_199# _336_/a_215_47# 0.03fF
C607 _458_/X _421_/X 0.01fF
C608 _487_/X VPWR 8.40fF
C609 _523_/X _504_/X 0.03fF
C610 _603_/Y _504_/X 0.79fF
C611 output19/a_27_47# _628_/Y 0.02fF
C612 _390_/D _559_/a_227_297# 0.03fF
C613 _503_/a_381_47# _473_/a_77_199# 0.04fF
C614 _519_/A _631_/A 0.67fF
C615 _420_/a_448_47# _420_/X 0.01fF
C616 _613_/X _633_/Y 0.43fF
C617 _457_/X _460_/a_226_47# 0.16fF
C618 _512_/a_78_199# _514_/A 0.21fF
C619 B[1] _330_/A 0.30fF
C620 _469_/a_62_47# _469_/a_381_47# 0.08fF
C621 _413_/X _561_/A 0.00fF
C622 _432_/A _432_/a_150_297# 0.03fF
C623 _630_/a_489_413# VPWR 0.41fF
C624 _566_/A _588_/A 0.26fF
C625 _380_/A _371_/B 0.03fF
C626 _625_/Y _610_/A 0.30fF
C627 _396_/a_250_297# _395_/X 0.18fF
C628 _387_/a_215_47# _350_/C 0.11fF
C629 _519_/a_183_297# VPWR 0.00fF
C630 _452_/A _418_/X 1.67fF
C631 _568_/a_323_297# _585_/B 0.04fF
C632 _540_/X _559_/a_77_199# 0.13fF
C633 VPWR _438_/X 1.34fF
C634 _634_/Y _442_/B 0.15fF
C635 _616_/Y _624_/a_76_199# 0.37fF
C636 _510_/X _511_/a_250_297# 0.20fF
C637 _381_/C VPWR 7.02fF
C638 _511_/a_93_21# _511_/a_250_297# 0.50fF
C639 _586_/a_76_199# _586_/a_218_47# 0.04fF
C640 M[1] _591_/A 0.19fF
C641 _465_/a_373_47# _464_/A 0.05fF
C642 _400_/a_80_21# _406_/A 0.20fF
C643 _507_/Y _483_/X 0.21fF
C644 _360_/a_489_413# _519_/A 0.09fF
C645 _548_/a_226_47# _530_/X 0.06fF
C646 _543_/Y _386_/A 0.39fF
C647 _607_/a_215_47# _601_/A 0.04fF
C648 _531_/B _531_/A 0.31fF
C649 _421_/a_226_47# VPWR 0.09fF
C650 _382_/B _383_/X 0.03fF
C651 _351_/a_27_53# B[5] 0.05fF
C652 _426_/A _397_/X 0.10fF
C653 _386_/A _515_/Y 0.35fF
C654 _616_/B _598_/A 0.73fF
C655 _440_/X _459_/a_226_47# 0.05fF
C656 _338_/X _337_/A 0.30fF
C657 _585_/B _584_/A 0.02fF
C658 _382_/B _356_/a_215_47# 0.16fF
C659 _410_/B _481_/A 0.03fF
C660 _538_/Y _485_/D 0.03fF
C661 B[0] _521_/a_215_47# 0.04fF
C662 _487_/X _559_/a_539_297# 0.02fF
C663 _459_/X _460_/a_226_47# 0.62fF
C664 input11/a_27_47# A[2] 0.01fF
C665 _402_/a_27_47# _433_/Y 0.14fF
C666 _492_/a_76_199# _492_/X 0.22fF
C667 _362_/a_489_413# _361_/X 0.14fF
C668 _569_/A _622_/C 0.04fF
C669 _410_/B _633_/Y 0.01fF
C670 _456_/a_226_47# _633_/Y 0.14fF
C671 _330_/A _383_/X 0.37fF
C672 VPWR _384_/a_76_199# 0.52fF
C673 _351_/X VPWR 1.66fF
C674 _628_/a_734_297# _621_/X 0.15fF
C675 VPWR _570_/A 3.51fF
C676 M[8] _464_/Y 0.01fF
C677 _375_/a_79_199# VPWR 0.64fF
C678 _443_/a_68_297# _443_/a_150_297# 0.02fF
C679 _571_/a_250_297# _570_/a_68_297# 0.03fF
C680 _595_/a_227_47# _595_/X 0.04fF
C681 _547_/X _515_/A 0.15fF
C682 _386_/a_664_47# _520_/X 0.08fF
C683 _502_/a_215_47# _527_/A 0.01fF
C684 VPWR _508_/a_77_199# 0.95fF
C685 VPWR _316_/a_62_47# 0.58fF
C686 _580_/A _576_/X 0.01fF
C687 _583_/X _607_/a_78_199# 0.05fF
C688 _503_/a_381_47# _471_/A 0.10fF
C689 _542_/C VPWR 5.13fF
C690 _555_/a_27_413# _555_/a_298_297# 0.02fF
C691 _375_/X _423_/a_78_199# 0.01fF
C692 _469_/a_558_47# _469_/X 0.24fF
C693 _538_/Y _483_/X 0.02fF
C694 _497_/B _462_/X 0.16fF
C695 _635_/a_27_413# _370_/B 0.03fF
C696 A[6] _507_/Y 0.08fF
C697 _365_/a_81_21# _371_/A 0.24fF
C698 _521_/X _521_/a_78_199# 0.21fF
C699 _582_/Y _602_/Y 0.00fF
C700 _567_/B _457_/X 0.77fF
C701 _445_/A _335_/a_381_47# 0.02fF
C702 VPWR _552_/a_226_47# 0.09fF
C703 _444_/Y _389_/a_27_47# 0.07fF
C704 _634_/Y _634_/a_27_413# 0.37fF
C705 _376_/X _481_/A 0.04fF
C706 _583_/X _591_/A 0.01fF
C707 _567_/B _467_/Y 0.03fF
C708 _475_/A _326_/A 0.61fF
C709 VPWR _430_/a_68_297# 0.27fF
C710 _554_/X VPWR 2.78fF
C711 _547_/X _535_/Y 0.09fF
C712 _627_/D _622_/C 0.33fF
C713 _406_/A _433_/Y 0.81fF
C714 _537_/a_77_199# _540_/a_93_21# 0.02fF
C715 _564_/a_219_297# _572_/A 0.17fF
C716 _621_/X _627_/B 2.02fF
C717 _485_/D _486_/X 0.11fF
C718 VPWR _535_/A 1.81fF
C719 _484_/a_78_199# _367_/C 0.01fF
C720 _352_/a_222_93# _328_/X 0.12fF
C721 _455_/X _587_/A 0.12fF
C722 A[5] VPWR 0.53fF
C723 _628_/a_382_297# _623_/a_489_413# 0.01fF
C724 _392_/A _631_/B 1.18fF
C725 _513_/A _485_/D 0.41fF
C726 M[2] _417_/A 1.17fF
C727 _587_/A _509_/A 0.42fF
C728 _412_/a_226_47# _631_/B 0.05fF
C729 _458_/X _460_/X 0.09fF
C730 _386_/X _515_/Y 1.40fF
C731 _635_/a_27_413# _371_/B 0.21fF
C732 _569_/Y _570_/X 0.37fF
C733 B[1] _442_/B 0.03fF
C734 _559_/X _588_/A 0.27fF
C735 _567_/B _459_/X 0.58fF
C736 _419_/X VPWR 12.14fF
C737 _485_/D _486_/a_150_297# 0.02fF
C738 _483_/X _486_/X 0.56fF
C739 _634_/a_300_297# VPWR 0.56fF
C740 _413_/X VPWR 1.21fF
C741 _563_/B _584_/A 0.21fF
C742 _439_/X _433_/Y 0.00fF
C743 _380_/A _361_/a_76_199# 0.02fF
C744 _583_/a_489_413# _602_/A 0.07fF
C745 _628_/a_300_47# _564_/a_27_53# 0.03fF
C746 _543_/A _503_/A 0.31fF
C747 _417_/D _417_/A 0.10fF
C748 input3/a_558_47# input3/a_664_47# 0.60fF
C749 input3/a_381_47# input3/a_841_47# 0.03fF
C750 _567_/B _503_/A 0.08fF
C751 _566_/A _559_/X 0.02fF
C752 _563_/A _519_/C 0.17fF
C753 _355_/a_161_47# _322_/A 0.04fF
C754 _497_/A VPWR 1.87fF
C755 B[7] _621_/X 0.35fF
C756 _516_/A _448_/B 0.83fF
C757 _359_/a_68_297# _359_/X 0.27fF
C758 _580_/A _549_/X 0.13fF
C759 _626_/Y output22/a_27_47# 0.60fF
C760 _557_/Y _558_/a_77_199# 0.37fF
C761 _623_/a_226_47# _627_/B 0.02fF
C762 _412_/a_226_47# _411_/X 0.57fF
C763 _417_/A _332_/X 0.03fF
C764 _386_/a_62_47# _386_/a_381_47# 0.08fF
C765 _444_/Y _411_/a_68_297# 0.01fF
C766 _456_/X _446_/X 2.87fF
C767 VPWR _629_/a_68_297# 0.27fF
C768 _442_/D _572_/A 0.28fF
C769 _457_/a_489_413# _504_/X 0.11fF
C770 _467_/Y _558_/a_77_199# 0.01fF
C771 _544_/A _379_/a_215_47# 0.05fF
C772 _491_/a_76_199# _491_/a_226_47# 0.49fF
C773 _594_/a_27_297# _573_/A 0.37fF
C774 _588_/Y _616_/A 0.09fF
C775 _448_/A _447_/B 0.16fF
C776 _315_/a_161_47# _449_/A 0.01fF
C777 _398_/a_226_297# _374_/X 0.02fF
C778 B[7] _624_/a_585_369# 0.01fF
C779 _633_/a_74_47# _633_/a_265_297# 0.03fF
C780 _524_/a_78_199# _525_/a_76_199# 0.02fF
C781 _419_/X _314_/X 0.12fF
C782 _490_/X _455_/X 0.02fF
C783 _623_/X _628_/Y 0.28fF
C784 output23/a_27_47# M[15] 0.44fF
C785 _588_/A _571_/a_93_21# 0.01fF
C786 _550_/a_78_199# _522_/a_226_47# 0.00fF
C787 A[6] _486_/X 0.16fF
C788 _429_/a_76_199# _398_/X 0.22fF
C789 _511_/a_250_297# _511_/X 0.03fF
C790 _446_/X _478_/A 0.03fF
C791 _429_/a_226_47# _397_/X 0.15fF
C792 _360_/a_76_199# _359_/X 0.29fF
C793 _370_/A B[5] 0.34fF
C794 _383_/X _442_/B 0.03fF
C795 _626_/a_109_297# _616_/A 0.02fF
C796 _626_/a_109_47# _616_/B 0.13fF
C797 _526_/a_76_199# _524_/X 0.02fF
C798 _526_/a_489_413# _504_/X 0.18fF
C799 _526_/a_226_47# _525_/X 0.53fF
C800 _463_/a_226_47# _464_/A 0.17fF
C801 _627_/A _539_/X 0.19fF
C802 _566_/A _571_/a_93_21# 0.20fF
C803 _533_/X _522_/a_226_47# 0.16fF
C804 _503_/a_62_47# _587_/A 0.10fF
C805 _597_/a_78_199# _597_/a_292_297# 0.03fF
C806 _513_/A A[6] 0.16fF
C807 _442_/D _620_/a_226_47# 0.00fF
C808 B[3] _620_/a_489_413# 0.01fF
C809 input12/a_381_47# _618_/Y 0.01fF
C810 _628_/a_300_47# _584_/A 0.45fF
C811 _569_/A _587_/A 0.24fF
C812 _485_/A _547_/a_222_93# 0.00fF
C813 _350_/C _332_/a_150_297# 0.01fF
C814 _422_/a_489_413# VPWR 0.39fF
C815 _569_/A _612_/A 0.21fF
C816 _512_/a_78_199# _512_/a_215_47# 0.26fF
C817 _423_/a_215_47# _396_/X 0.09fF
C818 _433_/Y _442_/A 0.16fF
C819 _498_/A _531_/A 0.30fF
C820 _350_/a_27_297# _350_/B 0.41fF
C821 _442_/D _542_/D 0.03fF
C822 output27/a_27_47# _432_/X 0.12fF
C823 _477_/a_493_297# VPWR 0.01fF
C824 _417_/D _484_/a_215_47# 0.16fF
C825 _371_/a_68_297# _432_/B 0.02fF
C826 _525_/a_489_413# VPWR 0.39fF
C827 _384_/X _397_/a_226_47# 0.33fF
C828 _506_/A _480_/A 0.08fF
C829 _539_/a_68_297# _587_/A 0.45fF
C830 _408_/X _408_/a_68_297# 0.27fF
C831 _390_/B _326_/A 0.03fF
C832 _586_/a_76_199# B[7] 0.10fF
C833 _627_/C _564_/a_27_53# 0.12fF
C834 _474_/A _533_/a_227_47# 0.02fF
C835 _497_/B _463_/a_76_199# 0.04fF
C836 _532_/a_76_199# _530_/X 0.12fF
C837 _576_/a_226_47# VPWR 0.18fF
C838 A[4] _390_/B 0.24fF
C839 _584_/A _322_/a_27_47# 0.02fF
C840 _336_/a_493_297# VPWR 0.01fF
C841 A[6] _454_/X 0.09fF
C842 _417_/D _469_/X 0.08fF
C843 _614_/a_76_199# _616_/A 0.22fF
C844 _567_/B _471_/Y 0.02fF
C845 _569_/A _625_/Y 0.07fF
C846 _386_/a_841_47# _386_/X 0.03fF
C847 A[3] _547_/X 0.03fF
C848 _590_/A _622_/X 0.45fF
C849 _588_/A _592_/a_113_297# 0.05fF
C850 _587_/A _627_/D 0.16fF
C851 _627_/D _612_/A 0.12fF
C852 _520_/X _537_/a_227_297# 0.03fF
C853 _428_/a_299_297# _428_/X 0.03fF
C854 _544_/A _567_/B 0.25fF
C855 _626_/Y _594_/X 0.07fF
C856 _585_/B _609_/a_80_21# 0.01fF
C857 _382_/a_68_297# _383_/a_489_413# 0.00fF
C858 _392_/Y _631_/B 0.56fF
C859 _494_/a_76_199# _494_/a_226_297# 0.01fF
C860 _494_/a_226_47# _494_/a_489_413# 0.02fF
C861 VPWR _489_/a_489_413# 0.39fF
C862 _366_/a_76_199# _366_/a_226_297# 0.01fF
C863 _366_/a_226_47# _366_/a_489_413# 0.02fF
C864 _487_/a_215_47# _487_/X 0.01fF
C865 VPWR _607_/a_292_297# 0.02fF
C866 _487_/X _563_/A 2.49fF
C867 _378_/a_664_47# _324_/a_558_47# 0.04fF
C868 _485_/A _518_/X 0.32fF
C869 _327_/a_292_297# _631_/A 0.02fF
C870 _314_/a_68_297# _328_/a_68_297# 0.01fF
C871 _608_/X _584_/A 0.02fF
C872 A[5] _399_/a_215_47# 0.33fF
C873 _461_/a_78_199# _422_/X 0.01fF
C874 _417_/D _512_/a_78_199# 0.12fF
C875 A[3] _570_/a_68_297# 0.03fF
C876 VPWR _540_/a_93_21# 0.40fF
C877 _338_/X VPWR 2.63fF
C878 _544_/A _565_/a_209_47# 0.03fF
C879 _471_/Y _468_/a_78_199# 0.01fF
C880 _550_/a_78_199# _521_/X 0.15fF
C881 _614_/a_489_413# M[1] 0.02fF
C882 VPWR _547_/a_544_297# 0.01fF
C883 _442_/D _478_/A 0.63fF
C884 _610_/A _433_/Y 0.02fF
C885 _596_/a_76_199# _626_/Y 0.08fF
C886 _575_/a_215_47# _548_/X 0.05fF
C887 _575_/a_493_297# _547_/X 0.08fF
C888 _353_/X _359_/X 1.47fF
C889 _324_/a_381_47# _367_/C 0.67fF
C890 _442_/a_27_47# _442_/A 0.48fF
C891 _599_/A _607_/a_78_199# 0.00fF
C892 _487_/X _627_/A 0.18fF
C893 _337_/A _631_/A 0.44fF
C894 _390_/D _328_/A 0.05fF
C895 VPWR _621_/X 2.18fF
C896 _347_/A _512_/a_78_199# 0.54fF
C897 _625_/Y _627_/D 0.28fF
C898 _533_/X _521_/X 0.51fF
C899 _597_/a_215_47# _574_/X 0.11fF
C900 _627_/C _584_/A 1.37fF
C901 VPWR _398_/X 1.19fF
C902 _586_/a_439_47# _503_/A 0.06fF
C903 _335_/a_62_47# VPWR 0.54fF
C904 _442_/D _619_/Y 0.00fF
C905 _567_/B _504_/X 0.03fF
C906 _513_/a_27_47# _542_/D 0.00fF
C907 _440_/a_489_413# _468_/X 0.01fF
C908 _464_/A _498_/A 0.02fF
C909 _413_/a_68_297# M[9] 0.01fF
C910 _381_/C _563_/A 1.39fF
C911 _432_/B _432_/X 0.01fF
C912 _445_/A _475_/A 2.03fF
C913 _451_/a_27_47# _451_/A 0.31fF
C914 input5/a_558_47# _478_/A 0.35fF
C915 _340_/A _530_/X 0.05fF
C916 _378_/A _367_/C 0.06fF
C917 _567_/B _566_/Y 0.31fF
C918 _551_/a_76_199# _552_/a_76_199# 0.05fF
C919 _627_/A _438_/X 0.28fF
C920 _332_/X _366_/a_76_199# 0.42fF
C921 _542_/A _472_/B 0.05fF
C922 _513_/A _418_/B 0.02fF
C923 _420_/X _391_/B 0.30fF
C924 _438_/a_68_297# _438_/X 0.27fF
C925 _532_/a_76_199# _557_/B 0.23fF
C926 _475_/A _350_/B 0.15fF
C927 _623_/X _624_/a_489_47# 0.01fF
C928 _346_/a_161_47# _442_/A 0.17fF
C929 _611_/X _616_/A 0.03fF
C930 _588_/A _530_/X 0.03fF
C931 _561_/A _485_/D 0.78fF
C932 _576_/X _616_/A 0.07fF
C933 _559_/X _616_/B 0.16fF
C934 _396_/a_250_297# _391_/A 0.00fF
C935 _315_/a_161_47# _417_/D 0.58fF
C936 _489_/a_226_47# _489_/a_76_199# 0.49fF
C937 _404_/a_664_47# _404_/a_841_47# 0.29fF
C938 _563_/A _570_/A 0.38fF
C939 _390_/D _389_/a_27_47# 0.23fF
C940 _347_/a_27_47# _417_/D 0.31fF
C941 _566_/A _530_/X 0.35fF
C942 _494_/a_489_413# _493_/X 0.14fF
C943 _623_/a_226_47# VPWR 0.08fF
C944 B[7] _485_/D 0.04fF
C945 output25/a_27_47# _351_/X 0.18fF
C946 _350_/X _398_/a_226_47# 0.01fF
C947 _366_/a_489_413# _337_/X 0.14fF
C948 _516_/A _514_/B 0.05fF
C949 _391_/B _411_/A 0.03fF
C950 _618_/A _625_/a_27_47# 0.17fF
C951 _461_/X _462_/a_76_199# 0.22fF
C952 _462_/X _462_/a_226_47# 0.05fF
C953 _347_/a_27_47# _347_/A 0.47fF
C954 _610_/A _610_/Y 1.68fF
C955 _627_/A _570_/A 0.53fF
C956 _356_/a_292_297# _452_/A 0.02fF
C957 _586_/a_76_199# VPWR 0.28fF
C958 B[1] _397_/X 0.01fF
C959 _586_/a_218_374# _622_/C 0.02fF
C960 _583_/X _557_/Y 0.01fF
C961 _602_/A _553_/a_78_199# 0.02fF
C962 input12/a_62_47# VPWR 0.53fF
C963 _443_/B _442_/A 0.10fF
C964 _456_/a_226_297# _454_/X 0.02fF
C965 _410_/B _334_/a_197_47# 0.07fF
C966 _583_/X _602_/A 0.51fF
C967 _550_/a_215_47# _550_/a_78_199# 0.26fF
C968 _511_/X _522_/X 2.24fF
C969 _631_/B _332_/X 0.21fF
C970 _630_/a_226_47# _629_/X 0.59fF
C971 _616_/A _618_/A 0.19fF
C972 _458_/X _390_/B 0.03fF
C973 _422_/a_76_199# _412_/X 0.34fF
C974 _532_/a_489_47# VPWR 0.05fF
C975 _342_/X _338_/X 0.32fF
C976 _424_/a_76_199# _423_/X 0.29fF
C977 _424_/a_226_47# _424_/X 0.05fF
C978 _452_/a_68_297# _449_/A 0.01fF
C979 _493_/X _458_/X 0.02fF
C980 _473_/a_77_199# _473_/a_227_297# 0.13fF
C981 _551_/a_489_413# _554_/A 0.01fF
C982 _362_/a_226_47# _351_/X 0.25fF
C983 _527_/B VPWR 1.90fF
C984 _542_/B _547_/X 0.03fF
C985 _633_/Y _385_/a_664_47# 0.08fF
C986 _543_/a_109_297# VPWR 0.02fF
C987 _318_/a_27_47# _485_/A 0.26fF
C988 _426_/A _427_/A 0.16fF
C989 _568_/a_227_47# VPWR 0.05fF
C990 _351_/a_27_53# _351_/X 0.03fF
C991 _382_/A VPWR 0.61fF
C992 _451_/a_27_47# _627_/B 0.01fF
C993 _561_/a_27_47# _454_/X 0.01fF
C994 _543_/B _544_/a_62_47# 0.10fF
C995 _417_/D _488_/a_226_47# 0.09fF
C996 _563_/A _419_/X 0.13fF
C997 _601_/A _624_/X 0.11fF
C998 _396_/a_250_297# _330_/A 0.10fF
C999 _448_/A _448_/a_68_297# 0.32fF
C1000 _567_/B _474_/Y 0.02fF
C1001 _561_/A A[6] 0.38fF
C1002 _436_/A _408_/a_68_297# 0.07fF
C1003 _506_/Y _507_/Y 0.51fF
C1004 _380_/A _378_/A 1.53fF
C1005 _538_/A _587_/A 0.02fF
C1006 _602_/A _580_/a_68_297# 0.02fF
C1007 _587_/A _510_/X 1.02fF
C1008 _587_/A _511_/a_93_21# 0.12fF
C1009 _517_/X _381_/B 0.37fF
C1010 _620_/a_226_47# _618_/A 0.06fF
C1011 _530_/a_76_199# _530_/a_226_47# 0.49fF
C1012 _442_/a_197_47# _442_/B 0.03fF
C1013 _455_/X _433_/Y 0.03fF
C1014 _542_/a_197_47# _542_/B 0.12fF
C1015 _469_/A _520_/X 0.70fF
C1016 _445_/A _390_/B 0.03fF
C1017 B[7] A[6] 0.37fF
C1018 _437_/a_222_93# VPWR 0.07fF
C1019 _622_/a_29_53# _622_/a_183_297# 0.04fF
C1020 _433_/Y _509_/A 0.09fF
C1021 _545_/Y _544_/a_381_47# 0.00fF
C1022 _399_/a_215_47# _398_/X 0.05fF
C1023 _594_/X _593_/A 0.30fF
C1024 _595_/a_539_297# _503_/A 0.08fF
C1025 _351_/A _350_/C 0.22fF
C1026 _510_/A VPWR 5.22fF
C1027 _482_/a_68_297# _347_/A 0.14fF
C1028 _572_/A _627_/a_27_297# 0.01fF
C1029 _327_/a_78_199# _328_/B 0.25fF
C1030 _583_/X _606_/A 2.10fF
C1031 _570_/A _537_/a_227_47# 0.39fF
C1032 _451_/a_27_47# B[7] 0.07fF
C1033 _391_/A _633_/Y 0.09fF
C1034 _627_/X _572_/A 0.14fF
C1035 _626_/Y _522_/a_76_199# 0.05fF
C1036 _331_/a_27_47# _383_/X 0.00fF
C1037 _418_/A _418_/X 1.15fF
C1038 _630_/a_226_47# _432_/B 0.25fF
C1039 _533_/X _580_/B 0.01fF
C1040 _551_/X _549_/X 0.23fF
C1041 _473_/a_323_297# _472_/Y 0.03fF
C1042 _626_/Y _492_/a_76_199# 0.02fF
C1043 _523_/a_76_199# _523_/a_226_297# 0.01fF
C1044 _523_/a_226_47# _523_/a_489_413# 0.02fF
C1045 VPWR _485_/D 4.47fF
C1046 _559_/X _530_/X 0.15fF
C1047 _363_/A B[5] 0.25fF
C1048 _587_/A _475_/A 0.23fF
C1049 _368_/a_68_297# _634_/a_27_413# 0.02fF
C1050 _608_/X _609_/a_80_21# 0.30fF
C1051 output27/a_27_47# M[4] 0.43fF
C1052 _447_/X M[9] 0.04fF
C1053 _456_/a_76_199# _456_/X 0.39fF
C1054 _532_/a_206_369# _527_/A 0.16fF
C1055 _532_/a_585_369# _527_/Y 0.05fF
C1056 _390_/D _631_/Y 0.08fF
C1057 _542_/D _627_/a_27_297# 0.25fF
C1058 B[7] _598_/B 0.06fF
C1059 _326_/a_27_47# _475_/A 0.07fF
C1060 _375_/a_222_93# _375_/a_448_47# 0.03fF
C1061 _352_/a_544_297# VPWR 0.01fF
C1062 _475_/X _503_/A 0.11fF
C1063 _455_/X _442_/a_27_47# 0.02fF
C1064 _396_/X _330_/A 0.03fF
C1065 _634_/a_300_297# _368_/A 0.12fF
C1066 _627_/C _609_/a_80_21# 0.00fF
C1067 _441_/a_292_297# _454_/X 0.02fF
C1068 _316_/a_381_47# _316_/a_664_47# 0.09fF
C1069 _548_/a_226_297# _546_/X 0.02fF
C1070 _538_/Y _559_/a_77_199# 0.41fF
C1071 _627_/X _542_/D 0.39fF
C1072 _476_/a_93_21# _471_/Y 0.08fF
C1073 _506_/A _585_/B 0.12fF
C1074 _508_/a_77_199# _508_/a_227_47# 0.24fF
C1075 VPWR _483_/X 2.62fF
C1076 _543_/Y _515_/A 0.03fF
C1077 _619_/Y _618_/A 1.04fF
C1078 output30/a_27_47# _557_/B 0.29fF
C1079 _537_/a_227_47# _535_/A 0.16fF
C1080 _530_/a_76_199# _529_/Y 0.22fF
C1081 _563_/D _547_/X 0.03fF
C1082 _566_/A _514_/B 0.25fF
C1083 _382_/B _481_/A 0.24fF
C1084 _580_/a_68_297# _606_/A 0.03fF
C1085 _515_/Y _515_/A 1.50fF
C1086 _485_/a_27_47# _563_/B 0.01fF
C1087 _595_/a_77_199# _595_/a_227_297# 0.13fF
C1088 VPWR _631_/A 7.74fF
C1089 _503_/a_62_47# _433_/Y 0.12fF
C1090 _569_/A _433_/Y 0.10fF
C1091 B[0] _514_/A 0.13fF
C1092 _536_/Y _472_/B 0.06fF
C1093 _561_/A _418_/B 0.62fF
C1094 _543_/Y _546_/a_76_199# 0.39fF
C1095 _410_/B _509_/Y 0.60fF
C1096 _515_/Y _546_/a_76_199# 0.00fF
C1097 _442_/D _381_/B 0.05fF
C1098 _516_/A _517_/a_68_297# 0.05fF
C1099 _440_/X _460_/a_226_297# 0.01fF
C1100 _455_/X _346_/a_161_47# 0.20fF
C1101 _574_/X _574_/a_299_297# 0.03fF
C1102 _604_/X _582_/a_27_47# 0.01fF
C1103 _608_/a_215_47# _608_/X 0.01fF
C1104 B[7] _549_/a_226_47# 0.06fF
C1105 _417_/D output29/a_27_47# 0.00fF
C1106 _359_/A _519_/A 0.76fF
C1107 _433_/Y _540_/a_250_297# 0.02fF
C1108 _554_/X _523_/X 0.19fF
C1109 _349_/a_215_47# _408_/B 0.16fF
C1110 _360_/a_489_413# VPWR 0.38fF
C1111 A[6] VPWR 3.35fF
C1112 _413_/X _419_/a_489_413# 0.07fF
C1113 _610_/A _621_/a_493_297# 0.08fF
C1114 _554_/X _603_/Y 0.42fF
C1115 _550_/X _530_/X 0.09fF
C1116 _627_/D _433_/Y 0.60fF
C1117 _559_/a_77_199# _486_/X 0.01fF
C1118 _556_/Y _558_/a_539_297# 0.04fF
C1119 _436_/A _436_/X 0.03fF
C1120 _455_/a_79_199# _413_/X 0.01fF
C1121 _494_/a_76_199# VPWR 0.50fF
C1122 _608_/a_215_47# _627_/C 0.20fF
C1123 _461_/a_215_47# VPWR 0.05fF
C1124 _498_/Y _527_/A 0.54fF
C1125 _410_/C _469_/X 0.25fF
C1126 _491_/a_226_47# _491_/X 0.05fF
C1127 _491_/a_76_199# _490_/X 0.32fF
C1128 _586_/S _627_/D 0.23fF
C1129 _506_/Y _454_/X 0.15fF
C1130 _539_/a_68_297# _540_/X 0.01fF
C1131 _410_/a_27_47# _442_/D 0.01fF
C1132 _633_/Y _632_/a_78_199# 0.01fF
C1133 _627_/C _627_/a_109_297# 0.04fF
C1134 _553_/a_78_199# _504_/X 0.33fF
C1135 _544_/A output32/a_27_47# 0.10fF
C1136 _455_/X _443_/B 0.15fF
C1137 _351_/A _380_/A 0.93fF
C1138 _423_/a_215_47# _423_/X 0.01fF
C1139 _416_/a_215_47# _418_/X 0.08fF
C1140 _458_/X _439_/a_226_47# 0.07fF
C1141 _452_/A _324_/a_381_47# 0.05fF
C1142 _451_/a_27_47# VPWR 0.54fF
C1143 _475_/X _471_/Y 0.36fF
C1144 _453_/X _453_/a_250_297# 0.03fF
C1145 _561_/a_27_47# _561_/A 0.31fF
C1146 _495_/a_76_199# _468_/X 0.42fF
C1147 _569_/Y _610_/A 0.03fF
C1148 B[4] _374_/a_78_199# 0.01fF
C1149 _519_/A _350_/C 0.09fF
C1150 _540_/X _540_/a_250_297# 0.03fF
C1151 _595_/a_539_297# _566_/Y 0.02fF
C1152 _412_/a_226_47# _408_/X 0.26fF
C1153 _338_/a_448_47# _332_/X 0.14fF
C1154 _534_/a_80_21# _530_/X 0.10fF
C1155 _547_/a_222_93# _547_/X 0.05fF
C1156 _425_/a_226_47# _426_/B 0.05fF
C1157 _383_/X _384_/a_489_413# 0.14fF
C1158 _612_/Y _624_/a_489_47# 0.13fF
C1159 _356_/a_78_199# _447_/B 0.05fF
C1160 _513_/a_27_47# _381_/B 0.00fF
C1161 B[6] VPWR 0.36fF
C1162 VPWR _391_/a_68_297# 0.32fF
C1163 _587_/A _390_/B 1.23fF
C1164 _349_/a_78_199# _419_/X 0.12fF
C1165 _378_/A _452_/A 0.51fF
C1166 _443_/A VPWR 1.27fF
C1167 _432_/A _371_/B 0.14fF
C1168 _587_/A _601_/A 0.01fF
C1169 input16/a_27_47# B[7] 0.45fF
C1170 _543_/Y _469_/a_664_47# 0.02fF
C1171 _598_/B VPWR 1.98fF
C1172 _342_/X _631_/A 0.03fF
C1173 _585_/B _535_/Y 0.13fF
C1174 _519_/A _367_/C 1.38fF
C1175 _623_/a_489_413# _433_/Y 0.11fF
C1176 _386_/a_841_47# _515_/A 0.05fF
C1177 _631_/Y _316_/a_558_47# 0.08fF
C1178 _578_/a_292_297# VPWR 0.01fF
C1179 _426_/B VPWR 1.10fF
C1180 _469_/A _503_/A 2.42fF
C1181 _482_/a_68_297# _477_/a_78_199# 0.01fF
C1182 _356_/a_78_199# _376_/a_68_297# 0.00fF
C1183 _340_/a_27_47# _445_/a_68_297# 0.00fF
C1184 _610_/Y _627_/D 0.05fF
C1185 _615_/a_215_47# _593_/Y 0.10fF
C1186 _475_/X _504_/X 0.00fF
C1187 _548_/a_76_199# _548_/a_226_297# 0.01fF
C1188 _548_/a_226_47# _548_/a_489_413# 0.02fF
C1189 _542_/B _480_/A 0.11fF
C1190 _359_/a_150_297# _383_/X 0.02fF
C1191 _436_/X _478_/A 0.27fF
C1192 _416_/a_493_297# _561_/A 0.02fF
C1193 _442_/D _542_/A 0.58fF
C1194 _584_/A _469_/X 0.60fF
C1195 _350_/a_205_297# _350_/C 0.02fF
C1196 _544_/A _485_/A 0.03fF
C1197 _393_/A _475_/A 0.32fF
C1198 _634_/a_300_297# _370_/A 0.00fF
C1199 _625_/Y _601_/A 0.24fF
C1200 _598_/a_68_297# _593_/Y 0.01fF
C1201 _628_/a_382_297# _623_/X 0.09fF
C1202 _360_/X _342_/a_68_297# 0.20fF
C1203 _516_/a_27_47# _570_/A 0.29fF
C1204 _599_/A _606_/A 0.13fF
C1205 _586_/S _541_/a_78_199# 0.01fF
C1206 _418_/B VPWR 1.27fF
C1207 _601_/Y _601_/A 0.38fF
C1208 _626_/Y _466_/X 0.35fF
C1209 _358_/a_27_47# _381_/B 0.30fF
C1210 _474_/A _476_/a_256_47# 0.02fF
C1211 _474_/Y _476_/a_93_21# 0.46fF
C1212 _542_/B _481_/A 0.15fF
C1213 _549_/a_226_47# VPWR 0.10fF
C1214 _337_/B _337_/X 0.01fF
C1215 _453_/a_250_297# _542_/D 0.03fF
C1216 _525_/a_489_413# _523_/X 0.07fF
C1217 _503_/A _559_/a_227_47# 0.50fF
C1218 _633_/Y _442_/B 0.05fF
C1219 _424_/a_489_413# VPWR 0.33fF
C1220 _469_/A _549_/a_76_199# 0.02fF
C1221 _442_/A _507_/Y 1.16fF
C1222 _587_/A _471_/A 0.58fF
C1223 _613_/a_227_47# _588_/A 0.02fF
C1224 _475_/a_68_297# _438_/X 0.01fF
C1225 _465_/X _467_/a_109_297# 0.01fF
C1226 _466_/X _467_/a_109_47# 0.67fF
C1227 _572_/B _571_/a_250_297# 0.03fF
C1228 _542_/C _478_/a_27_47# 0.30fF
C1229 _623_/X _622_/C 0.03fF
C1230 _387_/a_78_199# _409_/a_78_199# 0.03fF
C1231 _542_/A _521_/a_215_47# 0.02fF
C1232 _472_/Y VPWR 1.99fF
C1233 _539_/A _472_/B 1.52fF
C1234 _474_/A _478_/A 0.33fF
C1235 _563_/A _510_/A 0.05fF
C1236 B[7] _590_/B 0.08fF
C1237 _568_/a_323_297# _546_/X 0.03fF
C1238 _513_/a_27_47# _542_/A 0.20fF
C1239 _561_/a_27_47# VPWR 0.54fF
C1240 _510_/X _433_/Y 0.23fF
C1241 _538_/A _433_/Y 0.28fF
C1242 _544_/A _544_/a_841_47# 0.05fF
C1243 _511_/a_93_21# _433_/Y 0.15fF
C1244 _459_/a_76_199# _457_/X 0.35fF
C1245 _510_/A _627_/A 1.15fF
C1246 input16/a_27_47# VPWR 0.54fF
C1247 _510_/A _438_/a_68_297# 0.07fF
C1248 _589_/a_226_47# _590_/B 0.05fF
C1249 _563_/A _485_/D 0.44fF
C1250 _530_/X _557_/B 0.11fF
C1251 VPWR _446_/a_250_297# 0.74fF
C1252 _404_/a_664_47# _442_/D 0.20fF
C1253 _359_/B _381_/B 0.13fF
C1254 _567_/B _487_/X 0.06fF
C1255 _542_/D _514_/A 0.31fF
C1256 _417_/D _479_/B 0.03fF
C1257 _474_/Y _475_/X 0.86fF
C1258 _604_/a_80_21# _604_/a_209_297# 0.16fF
C1259 _390_/D _326_/A 0.38fF
C1260 VPWR _525_/X 2.21fF
C1261 input7/a_27_47# _542_/A 0.22fF
C1262 _452_/X _628_/Y 0.12fF
C1263 _353_/X _417_/A 0.83fF
C1264 _386_/X _412_/X 0.47fF
C1265 _504_/a_77_199# _504_/a_227_297# 0.13fF
C1266 _627_/A _485_/D 0.03fF
C1267 _359_/A _454_/X 0.12fF
C1268 _538_/A _540_/X 0.29fF
C1269 _497_/B _498_/Y 0.06fF
C1270 _369_/a_76_199# B[5] 0.17fF
C1271 _570_/X VPWR 1.07fF
C1272 _534_/a_80_21# _514_/B 0.29fF
C1273 _585_/B A[3] 0.25fF
C1274 _447_/a_68_297# _447_/X 0.27fF
C1275 _338_/X _370_/A 0.23fF
C1276 _436_/A _392_/A 0.07fF
C1277 _469_/A _566_/Y 0.03fF
C1278 _567_/B _438_/X 0.18fF
C1279 _416_/a_493_297# VPWR 0.01fF
C1280 _437_/X _439_/a_226_297# 0.04fF
C1281 _556_/A _558_/a_77_199# 0.17fF
C1282 _397_/a_76_199# _397_/a_489_413# 0.12fF
C1283 _436_/A _412_/a_226_47# 0.06fF
C1284 _459_/a_76_199# _459_/X 0.26fF
C1285 _563_/D _481_/A 0.30fF
C1286 _504_/a_77_199# _587_/A 0.02fF
C1287 _485_/D _548_/X 0.34fF
C1288 _479_/a_68_297# _505_/a_80_21# 0.02fF
C1289 _453_/X _449_/A 0.65fF
C1290 B[0] _417_/D 5.52fF
C1291 _627_/A _483_/X 0.03fF
C1292 _563_/D _633_/Y 0.03fF
C1293 _513_/A _367_/C 0.18fF
C1294 _556_/Y _530_/X 0.14fF
C1295 _560_/a_27_47# _627_/B 0.22fF
C1296 _343_/a_226_297# _329_/X 0.02fF
C1297 _437_/X VPWR 2.44fF
C1298 _347_/A B[0] 0.18fF
C1299 _417_/D _521_/a_292_297# 0.02fF
C1300 _488_/a_76_199# _520_/X 0.04fF
C1301 _490_/X _524_/X 0.01fF
C1302 _513_/A _442_/A 0.78fF
C1303 _426_/A _430_/X 1.13fF
C1304 _438_/X _468_/a_78_199# 0.15fF
C1305 _441_/a_292_297# VPWR 0.01fF
C1306 _562_/a_292_297# _584_/A 0.01fF
C1307 _587_/A _439_/a_226_47# 0.06fF
C1308 _486_/A _486_/a_68_297# 0.32fF
C1309 _581_/B VPWR 1.49fF
C1310 _523_/a_226_47# _522_/a_76_199# 0.01fF
C1311 _523_/a_76_199# _522_/a_226_47# 0.01fF
C1312 _439_/a_76_199# _439_/a_226_297# 0.01fF
C1313 _439_/a_226_47# _439_/a_489_413# 0.02fF
C1314 _371_/A _371_/B 3.03fF
C1315 _629_/B _373_/Y 0.76fF
C1316 _567_/B _570_/A 0.00fF
C1317 _508_/a_227_297# _507_/Y 0.03fF
C1318 _503_/a_62_47# _503_/a_558_47# 0.03fF
C1319 _603_/a_109_297# _579_/X 0.06fF
C1320 _338_/a_222_93# _338_/X 0.05fF
C1321 _420_/X _421_/a_226_47# 0.59fF
C1322 _540_/X _488_/X 0.06fF
C1323 _454_/X _367_/C 0.05fF
C1324 _487_/a_215_47# A[6] 0.08fF
C1325 _474_/Y _504_/a_539_297# 0.08fF
C1326 _569_/A _569_/Y 2.77fF
C1327 _563_/A A[6] 0.85fF
C1328 _530_/X _514_/B 0.09fF
C1329 _534_/a_209_297# _381_/B 0.12fF
C1330 _586_/S _586_/a_218_374# 0.02fF
C1331 _542_/B _515_/Y 0.05fF
C1332 _461_/X _478_/A 0.03fF
C1333 _543_/Y _542_/B 0.30fF
C1334 _627_/D _621_/a_493_297# 0.02fF
C1335 _635_/Y A[0] 0.42fF
C1336 _611_/a_27_297# _610_/A 0.52fF
C1337 _537_/a_323_297# _535_/Y 0.03fF
C1338 _418_/a_68_297# _378_/a_381_47# 0.01fF
C1339 _454_/X _442_/A 1.10fF
C1340 _392_/A _350_/X 0.48fF
C1341 _376_/X _417_/A 0.03fF
C1342 VPWR _439_/a_76_199# 0.50fF
C1343 _629_/B VPWR 1.69fF
C1344 _455_/X _519_/A 0.65fF
C1345 _590_/B VPWR 2.06fF
C1346 _621_/a_215_47# _621_/X 0.01fF
C1347 _627_/A A[6] 0.16fF
C1348 _587_/A _573_/Y 0.21fF
C1349 _603_/Y _527_/B 0.08fF
C1350 _616_/A _593_/Y 0.03fF
C1351 _396_/X _397_/X 0.15fF
C1352 _594_/X _598_/A 0.07fF
C1353 _609_/a_80_21# _469_/X 0.21fF
C1354 _623_/X _612_/A 3.14fF
C1355 _563_/A _451_/a_27_47# 0.02fF
C1356 _386_/A _411_/X 0.01fF
C1357 _605_/a_209_297# VPWR 0.45fF
C1358 _633_/Y _489_/a_226_47# 0.14fF
C1359 _569_/Y _627_/D 0.22fF
C1360 _361_/a_226_47# _361_/a_489_413# 0.02fF
C1361 _634_/Y B[5] 0.54fF
C1362 input3/a_664_47# _616_/B 0.02fF
C1363 _328_/a_68_297# _328_/a_150_297# 0.02fF
C1364 _462_/a_226_47# _462_/a_489_413# 0.02fF
C1365 _462_/a_76_199# _462_/a_226_297# 0.01fF
C1366 M[8] _501_/a_109_47# 0.14fF
C1367 _596_/a_76_199# _598_/A 0.37fF
C1368 _544_/a_62_47# VPWR 0.64fF
C1369 _449_/A _542_/D 0.36fF
C1370 _544_/a_381_47# _544_/a_558_47# 0.32fF
C1371 _506_/Y VPWR 2.42fF
C1372 _630_/X _398_/a_226_47# 0.07fF
C1373 _556_/Y _557_/B 0.46fF
C1374 _410_/B _469_/X 0.34fF
C1375 _633_/Y _591_/A 1.37fF
C1376 _623_/X _625_/Y 2.26fF
C1377 M[8] VPWR 2.00fF
C1378 _443_/a_68_297# _443_/B 0.30fF
C1379 _478_/A _431_/X 0.03fF
C1380 _523_/a_76_199# _521_/X 0.01fF
C1381 _622_/C _469_/a_841_47# 0.06fF
C1382 _513_/A _380_/A 0.72fF
C1383 _509_/A _507_/Y 0.27fF
C1384 _337_/A _367_/C 1.06fF
C1385 _473_/a_77_199# _433_/Y 0.18fF
C1386 _476_/X VPWR 2.06fF
C1387 _567_/B _497_/A 0.05fF
C1388 _496_/a_78_199# VPWR 0.63fF
C1389 _619_/a_27_47# _599_/A 0.03fF
C1390 _486_/A _486_/B 1.31fF
C1391 _390_/B _433_/Y 0.27fF
C1392 _386_/X _631_/B 1.01fF
C1393 _404_/a_381_47# _503_/A 0.61fF
C1394 VPWR _559_/a_77_199# 0.91fF
C1395 _524_/a_215_47# _626_/Y 0.11fF
C1396 _388_/a_27_47# VPWR 0.53fF
C1397 _549_/X _551_/a_489_413# 0.07fF
C1398 _417_/A M[9] 0.18fF
C1399 _386_/A _505_/a_303_47# 0.05fF
C1400 _419_/X _420_/X 2.78fF
C1401 _612_/Y _624_/X 0.36fF
C1402 _516_/A _517_/X 0.18fF
C1403 M[13] _620_/X 0.30fF
C1404 _627_/A _609_/a_209_47# 0.01fF
C1405 _503_/A _547_/X 0.03fF
C1406 _380_/A _454_/X 0.03fF
C1407 _574_/X _547_/X 1.06fF
C1408 _386_/a_664_47# _570_/A 0.08fF
C1409 _433_/a_109_47# _431_/X 0.23fF
C1410 _335_/a_381_47# _335_/a_664_47# 0.09fF
C1411 _380_/A _334_/a_27_47# 0.02fF
C1412 _336_/a_215_47# _519_/A 0.27fF
C1413 _563_/D _515_/Y 0.10fF
C1414 _542_/C _386_/a_664_47# 0.19fF
C1415 _351_/X _374_/X 0.06fF
C1416 _386_/X _411_/X 0.25fF
C1417 VPWR _394_/a_664_47# 0.38fF
C1418 _503_/A _570_/a_68_297# 0.14fF
C1419 _390_/D _445_/A 0.10fF
C1420 _615_/a_215_47# _595_/X 0.05fF
C1421 M[8] _501_/Y 0.76fF
C1422 _448_/B _378_/a_62_47# 0.02fF
C1423 _491_/X _490_/X 0.45fF
C1424 _465_/a_109_297# VPWR 0.39fF
C1425 _448_/A _378_/A 0.02fF
C1426 _417_/D _418_/a_68_297# 0.15fF
C1427 _400_/a_209_47# _391_/B 0.01fF
C1428 _496_/a_78_199# _496_/a_215_47# 0.26fF
C1429 _478_/a_197_47# _410_/C 0.03fF
C1430 _560_/a_27_47# VPWR 0.54fF
C1431 _528_/a_81_21# VPWR 0.49fF
C1432 _595_/a_227_47# A[3] 0.11fF
C1433 A[6] _505_/a_209_297# 0.14fF
C1434 _454_/X _316_/a_381_47# 0.12fF
C1435 _559_/a_77_199# _559_/a_539_297# 0.06fF
C1436 _520_/X _480_/A 0.07fF
C1437 _612_/Y _622_/C 0.13fF
C1438 _411_/a_150_297# _475_/A 0.01fF
C1439 _631_/a_109_297# _631_/Y 0.02fF
C1440 _361_/a_226_47# _361_/a_76_199# 0.49fF
C1441 _485_/a_27_47# _484_/a_215_47# 0.04fF
C1442 B[1] B[5] 0.63fF
C1443 _546_/a_489_413# VPWR 0.39fF
C1444 _402_/a_27_47# VPWR 0.53fF
C1445 _471_/A _433_/Y 0.03fF
C1446 _610_/Y _601_/A 0.00fF
C1447 _387_/a_292_297# VPWR 0.01fF
C1448 _549_/a_489_413# _540_/X 0.07fF
C1449 _549_/a_226_47# _548_/X 0.51fF
C1450 _577_/a_226_47# _580_/A 0.05fF
C1451 _360_/X _408_/B 0.03fF
C1452 _511_/a_250_297# _631_/Y 0.21fF
C1453 _480_/Y _442_/D 0.03fF
C1454 _627_/A _472_/Y 0.05fF
C1455 _539_/a_68_297# _507_/Y 0.06fF
C1456 A[5] _374_/X 0.17fF
C1457 _561_/A _367_/C 0.07fF
C1458 _612_/Y _618_/Y 0.06fF
C1459 _596_/a_226_47# _599_/Y 0.00fF
C1460 _445_/A _328_/A 0.48fF
C1461 _467_/a_109_47# _467_/a_397_297# 0.05fF
C1462 _554_/A _554_/a_68_297# 0.32fF
C1463 VPWR _399_/a_78_199# 0.60fF
C1464 _515_/Y _518_/a_250_297# 0.03fF
C1465 _627_/C A[3] 0.03fF
C1466 _520_/X _481_/A 0.01fF
C1467 _513_/A _455_/X 0.15fF
C1468 _440_/X _493_/a_78_199# 0.33fF
C1469 _385_/a_62_47# _394_/a_62_47# 0.00fF
C1470 _465_/a_109_297# _501_/Y 0.12fF
C1471 _417_/D _542_/D 0.59fF
C1472 _436_/A _332_/X 0.01fF
C1473 _572_/a_68_297# _572_/a_150_297# 0.02fF
C1474 _520_/X _633_/Y 0.03fF
C1475 _532_/a_76_199# _532_/a_206_369# 0.69fF
C1476 _360_/X input6/a_27_47# 0.00fF
C1477 _329_/a_76_199# _329_/a_226_47# 0.49fF
C1478 _633_/Y _590_/A 0.03fF
C1479 _607_/X _442_/D 0.02fF
C1480 _516_/A _442_/D 0.03fF
C1481 _442_/D _539_/A 0.03fF
C1482 _544_/A _547_/X 0.24fF
C1483 _525_/a_76_199# _492_/X 0.01fF
C1484 _520_/a_76_199# _520_/a_489_413# 0.12fF
C1485 _383_/a_76_199# _383_/a_489_413# 0.12fF
C1486 _497_/a_68_297# VPWR 0.25fF
C1487 _406_/A VPWR 6.07fF
C1488 M[5] VPWR 1.07fF
C1489 _487_/X _537_/a_227_297# 0.01fF
C1490 _378_/A _418_/A 0.38fF
C1491 _406_/Y _461_/X 0.56fF
C1492 _317_/a_27_47# VPWR 0.66fF
C1493 _599_/Y _624_/a_76_199# 0.03fF
C1494 _452_/X _447_/B 0.00fF
C1495 _455_/X _454_/X 2.40fF
C1496 _409_/a_215_47# _445_/a_68_297# 0.03fF
C1497 _351_/A _475_/A 0.01fF
C1498 _338_/X _363_/A 0.01fF
C1499 _360_/X _375_/X 0.03fF
C1500 _460_/a_76_199# _460_/X 0.22fF
C1501 _338_/X _420_/X 0.18fF
C1502 _340_/A _517_/X 0.05fF
C1503 _479_/A _517_/X 0.00fF
C1504 _454_/X _509_/A 0.34fF
C1505 VPWR _428_/X 1.16fF
C1506 input13/a_27_47# _352_/X 0.02fF
C1507 _627_/A _570_/X 0.73fF
C1508 _610_/A _620_/X 0.08fF
C1509 _390_/B _443_/B 0.23fF
C1510 _426_/A _430_/a_68_297# 0.12fF
C1511 VPWR _531_/a_193_297# 0.01fF
C1512 M[2] _369_/a_489_413# 0.11fF
C1513 _538_/Y _540_/a_250_297# 0.18fF
C1514 _494_/a_226_47# _494_/X 0.05fF
C1515 _533_/X _552_/a_76_199# 0.38fF
C1516 _631_/B _395_/X 0.29fF
C1517 output22/a_27_47# _465_/X 0.01fF
C1518 _419_/a_76_199# _418_/X 0.22fF
C1519 _479_/B _410_/C 0.26fF
C1520 _385_/a_62_47# _385_/a_558_47# 0.03fF
C1521 input12/a_381_47# input12/a_664_47# 0.09fF
C1522 _359_/A VPWR 1.25fF
C1523 _455_/a_79_199# _418_/B 0.22fF
C1524 VPWR _555_/a_27_413# 0.38fF
C1525 _568_/a_77_199# _568_/a_227_297# 0.13fF
C1526 _396_/a_93_21# _391_/a_68_297# 0.01fF
C1527 M[13] VPWR 0.74fF
C1528 _439_/X VPWR 1.55fF
C1529 _379_/a_215_47# _382_/A 0.01fF
C1530 _566_/Y _547_/X 0.30fF
C1531 _347_/A _346_/A 0.72fF
C1532 B[7] _610_/A 2.01fF
C1533 _515_/Y _518_/X 0.04fF
C1534 _407_/a_27_47# _406_/Y 0.03fF
C1535 M[8] _531_/C 0.68fF
C1536 _322_/A _481_/A 0.99fF
C1537 _393_/A _394_/a_841_47# 0.34fF
C1538 _480_/A _483_/a_250_297# 0.08fF
C1539 _380_/A _561_/A 0.13fF
C1540 VPWR _350_/C 3.50fF
C1541 _532_/a_76_199# _498_/Y 0.03fF
C1542 _468_/X _458_/X 0.03fF
C1543 VPWR output26/a_27_47# 0.75fF
C1544 _338_/X _328_/X 0.02fF
C1545 _585_/B _591_/A 0.10fF
C1546 B[0] _410_/C 0.39fF
C1547 _378_/a_841_47# VPWR 0.39fF
C1548 _356_/a_78_199# _356_/a_292_297# 0.03fF
C1549 _563_/D _563_/B 0.08fF
C1550 _487_/a_78_199# VPWR 0.63fF
C1551 _422_/a_76_199# _422_/X 0.22fF
C1552 _440_/X _406_/Y 0.01fF
C1553 _390_/D _587_/A 0.10fF
C1554 _614_/a_489_413# _633_/Y 0.09fF
C1555 _567_/B _532_/a_489_47# 0.13fF
C1556 _612_/Y _612_/A 0.74fF
C1557 _471_/A _443_/B 0.00fF
C1558 VPWR _367_/C 5.53fF
C1559 _416_/a_215_47# _324_/a_381_47# 0.02fF
C1560 _469_/A _539_/X 0.27fF
C1561 _567_/B _527_/B 0.46fF
C1562 _350_/a_27_297# _350_/a_205_297# 0.01fF
C1563 _543_/a_109_297# _543_/A 0.01fF
C1564 _530_/a_226_47# _530_/X 0.05fF
C1565 _626_/Y _593_/Y 0.03fF
C1566 _513_/A _547_/a_448_47# 0.02fF
C1567 _493_/X _494_/X 0.71fF
C1568 VPWR _442_/A 8.15fF
C1569 B[3] _442_/D 0.07fF
C1570 A[2] VPWR 0.73fF
C1571 _623_/X _433_/Y 1.03fF
C1572 _568_/a_227_297# _566_/A 0.01fF
C1573 _335_/a_841_47# _631_/A 0.35fF
C1574 _399_/a_78_199# _399_/a_215_47# 0.26fF
C1575 _568_/a_227_47# _567_/B 0.11fF
C1576 _571_/a_250_297# _469_/X 0.03fF
C1577 _631_/Y _522_/X 0.14fF
C1578 _416_/a_215_47# _378_/A 0.13fF
C1579 _527_/A _531_/B 0.02fF
C1580 _616_/a_109_297# _616_/Y 0.02fF
C1581 _340_/A _442_/D 0.34fF
C1582 _625_/Y _612_/Y 3.76fF
C1583 _623_/X _586_/S 0.22fF
C1584 _580_/B M[0] 0.17fF
C1585 _374_/X _398_/X 0.55fF
C1586 _499_/a_299_297# VPWR 0.67fF
C1587 _542_/A _514_/A 0.18fF
C1588 _600_/a_27_297# _598_/B 0.48fF
C1589 _515_/Y _520_/X 0.06fF
C1590 _506_/Y _627_/A 0.20fF
C1591 _466_/a_215_47# _432_/X 0.07fF
C1592 _466_/a_493_297# _430_/X 0.12fF
C1593 _381_/C _485_/A 3.22fF
C1594 _594_/X _616_/B 0.26fF
C1595 _635_/Y _635_/a_300_297# 0.22fF
C1596 _628_/a_382_297# _628_/Y 0.29fF
C1597 _338_/X _329_/X 2.07fF
C1598 _442_/D _588_/A 0.06fF
C1599 _632_/a_493_297# VPWR 0.01fF
C1600 _559_/a_227_47# _539_/X 0.05fF
C1601 B[0] _584_/A 0.43fF
C1602 _607_/a_78_199# _616_/Y 0.13fF
C1603 M[5] _399_/a_215_47# 0.27fF
C1604 _463_/a_226_47# _406_/Y 0.25fF
C1605 _463_/a_76_199# _462_/X 0.22fF
C1606 _326_/a_27_47# _328_/A 0.02fF
C1607 _567_/B _510_/A 0.19fF
C1608 _566_/A _442_/D 0.03fF
C1609 _596_/a_76_199# _616_/B 0.05fF
C1610 _519_/A _475_/A 0.03fF
C1611 _595_/X _572_/A 0.03fF
C1612 _376_/X _382_/a_68_297# 0.00fF
C1613 input5/a_381_47# input5/a_558_47# 0.32fF
C1614 _577_/a_76_199# _559_/X 0.32fF
C1615 _627_/A _559_/a_77_199# 0.23fF
C1616 _337_/A _452_/A 0.06fF
C1617 _523_/X _525_/X 0.35fF
C1618 _535_/Y _469_/X 0.03fF
C1619 _603_/Y _525_/X 0.11fF
C1620 _503_/a_558_47# _473_/a_77_199# 0.01fF
C1621 _457_/X _460_/a_489_413# 0.00fF
C1622 _342_/X _350_/C 0.03fF
C1623 _588_/A _588_/Y 0.29fF
C1624 _610_/A VPWR 5.65fF
C1625 _633_/Y _503_/A 0.03fF
C1626 _487_/X _469_/A 0.75fF
C1627 _469_/a_62_47# _469_/a_558_47# 0.03fF
C1628 _386_/A _479_/B 0.42fF
C1629 _567_/B _485_/D 0.09fF
C1630 _479_/a_68_297# _486_/X 0.20fF
C1631 _623_/X _610_/Y 0.42fF
C1632 _396_/a_250_297# _391_/B 0.01fF
C1633 _417_/A _343_/a_489_413# 0.09fF
C1634 _634_/Y _351_/X 0.11fF
C1635 _513_/A _380_/a_27_47# 0.22fF
C1636 _529_/Y _530_/X 0.02fF
C1637 _540_/X _559_/a_227_297# 0.03fF
C1638 _386_/a_558_47# _479_/a_68_297# 0.01fF
C1639 _533_/X _489_/a_226_47# 0.05fF
C1640 _538_/A _538_/Y 1.51fF
C1641 _616_/Y _624_/a_206_369# 0.29fF
C1642 _616_/A _624_/a_76_199# 0.29fF
C1643 _511_/a_93_21# _511_/a_256_47# 0.03fF
C1644 _607_/X _618_/A 0.05fF
C1645 _437_/a_222_93# _411_/A 0.01fF
C1646 _380_/A VPWR 7.19fF
C1647 _520_/a_226_297# A[6] 0.02fF
C1648 _400_/a_209_297# _406_/A 0.04fF
C1649 _548_/a_489_413# _530_/X 0.11fF
C1650 _426_/A _398_/X 0.12fF
C1651 _382_/B _417_/A 0.99fF
C1652 _510_/A _411_/A 0.26fF
C1653 _421_/a_489_413# VPWR 0.39fF
C1654 _567_/B _483_/X 1.04fF
C1655 _520_/X _585_/B 0.41fF
C1656 _351_/a_301_297# B[5] 0.01fF
C1657 _386_/A B[0] 0.25fF
C1658 _585_/B _590_/A 0.15fF
C1659 _380_/a_27_47# _334_/a_27_47# 0.00fF
C1660 _563_/D _627_/C 0.31fF
C1661 _459_/X _460_/a_489_413# 0.14fF
C1662 _571_/a_250_297# _546_/X 0.21fF
C1663 _492_/a_226_47# _492_/X 0.05fF
C1664 _603_/Y _581_/B 0.22fF
C1665 _513_/a_27_47# _566_/A 0.10fF
C1666 _408_/B _314_/a_68_297# 0.44fF
C1667 _417_/A _330_/A 0.03fF
C1668 _614_/a_76_199# _588_/A 0.03fF
C1669 _569_/Y _595_/a_77_199# 0.16fF
C1670 VPWR _384_/a_226_47# 0.09fF
C1671 _375_/a_222_93# VPWR 0.06fF
C1672 _402_/a_27_47# _438_/a_68_297# 0.02fF
C1673 VPWR _316_/a_381_47# 0.31fF
C1674 _469_/A _570_/A 0.45fF
C1675 _386_/a_841_47# _520_/X 0.14fF
C1676 B[0] _521_/X 0.18fF
C1677 VPWR _508_/a_227_297# 0.01fF
C1678 _577_/a_76_199# _550_/X 0.02fF
C1679 _503_/a_558_47# _471_/A 0.08fF
C1680 _555_/a_215_297# _555_/a_298_297# 0.18fF
C1681 _469_/a_664_47# _469_/X 0.12fF
C1682 _420_/X _631_/A 1.44fF
C1683 _497_/B _461_/X 0.01fF
C1684 _538_/Y _488_/X 0.01fF
C1685 _449_/A _542_/A 0.03fF
C1686 _538_/A _486_/X 0.02fF
C1687 _365_/a_81_21# _371_/B 0.08fF
C1688 _561_/A _452_/A 0.58fF
C1689 _365_/a_299_297# _371_/A 0.03fF
C1690 _635_/a_300_297# _370_/B 0.23fF
C1691 _557_/Y _602_/Y 0.20fF
C1692 _546_/a_76_199# _546_/X 0.22fF
C1693 _602_/A _602_/Y 0.36fF
C1694 _451_/A _541_/a_78_199# 0.06fF
C1695 _633_/Y _471_/Y 0.05fF
C1696 _567_/B A[6] 0.05fF
C1697 _544_/A _481_/A 0.14fF
C1698 _506_/Y _508_/a_227_47# 0.09fF
C1699 _634_/Y _634_/a_300_297# 0.22fF
C1700 VPWR _552_/a_489_413# 0.39fF
C1701 B[7] _452_/A 0.39fF
C1702 _374_/a_215_47# _361_/X 0.30fF
C1703 _583_/X _621_/X 0.61fF
C1704 _627_/D _627_/B 0.92fF
C1705 _447_/B _376_/a_68_297# 0.33fF
C1706 _406_/B _433_/Y 0.13fF
C1707 _398_/a_76_199# _398_/a_226_47# 0.49fF
C1708 _569_/A B[7] 0.30fF
C1709 _537_/a_77_199# _540_/a_250_297# 0.07fF
C1710 _564_/a_27_53# _572_/A 0.03fF
C1711 _621_/X _622_/X 2.16fF
C1712 _417_/D _381_/B 0.23fF
C1713 _627_/C _586_/a_505_21# 0.06fF
C1714 _520_/a_226_47# _486_/B 0.01fF
C1715 _593_/A _593_/Y 2.92fF
C1716 _484_/a_78_199# _486_/A 0.21fF
C1717 _352_/a_79_199# _352_/X 0.29fF
C1718 _628_/a_734_297# _623_/a_489_413# 0.02fF
C1719 _338_/X _369_/a_76_199# 0.01fF
C1720 _559_/a_227_47# _570_/A 0.10fF
C1721 _347_/A _381_/B 0.41fF
C1722 _444_/Y _443_/B 0.30fF
C1723 _468_/X _587_/A 0.07fF
C1724 _598_/a_68_297# _575_/X 0.00fF
C1725 _510_/X _454_/X 0.58fF
C1726 B[1] _384_/a_76_199# 0.05fF
C1727 _454_/X _511_/a_93_21# 0.07fF
C1728 _633_/Y _391_/B 0.03fF
C1729 _611_/X _588_/A 0.03fF
C1730 _633_/Y _504_/X 0.21fF
C1731 _386_/X B[0] 0.08fF
C1732 _567_/B B[6] 0.01fF
C1733 _627_/C _591_/A 1.52fF
C1734 _455_/X VPWR 6.60fF
C1735 _582_/a_27_47# _582_/Y 0.11fF
C1736 _582_/a_109_297# _557_/Y 0.06fF
C1737 _476_/X _523_/X 0.30fF
C1738 _583_/a_226_297# _602_/A 0.04fF
C1739 _488_/X _486_/X 0.84fF
C1740 A[3] _469_/X 0.70fF
C1741 B[7] _627_/D 1.43fF
C1742 input3/a_558_47# input3/a_841_47# 0.07fF
C1743 _381_/C _383_/X 0.02fF
C1744 _635_/a_27_413# VPWR 0.37fF
C1745 VPWR _509_/A 1.09fF
C1746 _580_/A _580_/B 0.86fF
C1747 B[0] _550_/a_215_47# 0.01fF
C1748 _412_/a_489_413# _411_/X 0.14fF
C1749 _563_/A _350_/C 0.41fF
C1750 _584_/A _572_/A 0.40fF
C1751 _623_/a_489_413# _627_/B 0.13fF
C1752 _386_/a_62_47# _386_/a_558_47# 0.03fF
C1753 _344_/a_78_199# _344_/a_215_47# 0.26fF
C1754 _623_/a_226_47# _622_/X 0.54fF
C1755 _520_/X _550_/a_78_199# 0.01fF
C1756 _587_/A _631_/Y 0.03fF
C1757 _512_/a_215_47# _542_/A 0.27fF
C1758 _420_/X _391_/a_68_297# 0.07fF
C1759 _391_/A _631_/B 0.03fF
C1760 _577_/a_76_199# _530_/X 0.10fF
C1761 _328_/B _519_/A 0.26fF
C1762 _457_/a_226_297# _504_/X 0.01fF
C1763 _491_/a_76_199# _491_/a_489_413# 0.12fF
C1764 _594_/a_109_297# _573_/A 0.12fF
C1765 _533_/X _520_/X 0.31fF
C1766 _611_/a_109_297# _591_/A 0.32fF
C1767 _487_/a_78_199# _487_/a_215_47# 0.26fF
C1768 _554_/a_68_297# _554_/a_150_297# 0.02fF
C1769 _602_/Y _606_/A 0.02fF
C1770 input8/a_27_47# VPWR 0.60fF
C1771 _436_/A _584_/A 0.82fF
C1772 _530_/a_76_199# _531_/B 0.32fF
C1773 _608_/a_78_199# _584_/A 0.28fF
C1774 _524_/a_78_199# _525_/a_226_47# 0.02fF
C1775 _478_/A _410_/C 0.47fF
C1776 _383_/X _384_/a_76_199# 0.27fF
C1777 _337_/a_68_297# _337_/a_150_297# 0.02fF
C1778 _550_/a_78_199# _522_/a_489_413# 0.01fF
C1779 _429_/a_226_47# _398_/X 0.55fF
C1780 _417_/A _442_/B 1.49fF
C1781 _313_/a_27_47# _395_/a_68_297# 0.00fF
C1782 _360_/a_226_47# _359_/X 0.53fF
C1783 VPWR _621_/a_78_199# 0.61fF
C1784 _563_/A _442_/A 0.40fF
C1785 _626_/a_397_297# _616_/A 0.14fF
C1786 _550_/X _522_/a_76_199# 0.01fF
C1787 _510_/a_68_297# _471_/Y 0.01fF
C1788 _527_/B _553_/a_78_199# 0.01fF
C1789 _526_/a_226_47# _524_/X 0.01fF
C1790 _526_/a_226_297# _504_/X 0.04fF
C1791 _526_/a_489_413# _525_/X 0.16fF
C1792 B[1] _419_/X 0.08fF
C1793 _584_/A _542_/D 0.13fF
C1794 _442_/D _620_/a_489_413# 0.00fF
C1795 _503_/a_381_47# _587_/A 0.12fF
C1796 _591_/Y _633_/Y 0.24fF
C1797 VPWR _397_/a_76_199# 0.57fF
C1798 _408_/B _313_/A 0.25fF
C1799 B[4] VPWR 0.54fF
C1800 _390_/D _433_/Y 0.12fF
C1801 _612_/Y _433_/Y 0.07fF
C1802 _393_/A _363_/a_68_297# 0.08fF
C1803 _477_/a_215_47# VPWR 0.06fF
C1804 _519_/a_29_53# _542_/A 0.37fF
C1805 _384_/X _397_/a_489_413# 0.07fF
C1806 _452_/A VPWR 3.67fF
C1807 _627_/A _442_/A 0.03fF
C1808 _539_/a_150_297# _587_/A 0.02fF
C1809 _417_/D _542_/A 1.16fF
C1810 _561_/A _541_/a_78_199# 0.01fF
C1811 _612_/Y _586_/S 0.26fF
C1812 _497_/B _463_/a_226_47# 0.13fF
C1813 _503_/a_62_47# VPWR 0.51fF
C1814 _576_/a_489_413# VPWR 0.43fF
C1815 _569_/A VPWR 2.24fF
C1816 _454_/a_556_47# _453_/X 0.02fF
C1817 _626_/Y _525_/a_76_199# 0.08fF
C1818 _585_/B _503_/A 0.20fF
C1819 _506_/Y _533_/a_323_297# 0.02fF
C1820 _347_/A _542_/A 0.16fF
C1821 _557_/Y _558_/X 0.04fF
C1822 _336_/a_215_47# VPWR 0.05fF
C1823 _614_/a_226_47# _616_/A 0.05fF
C1824 _441_/a_215_47# _355_/A 0.24fF
C1825 _569_/Y _623_/X 0.05fF
C1826 _584_/A _350_/X 0.15fF
C1827 _544_/A _543_/Y 1.01fF
C1828 _545_/Y _622_/C 0.81fF
C1829 A[3] _546_/X 0.03fF
C1830 _588_/A _592_/a_199_47# 0.05fF
C1831 _539_/X _570_/a_68_297# 0.02fF
C1832 _520_/X _537_/a_323_297# 0.03fF
C1833 _505_/a_209_47# _482_/X 0.01fF
C1834 _544_/A _515_/Y 0.02fF
C1835 _581_/a_27_93# _583_/a_76_199# 0.00fF
C1836 _539_/a_68_297# VPWR 0.32fF
C1837 _421_/X VPWR 1.27fF
C1838 _390_/D _540_/X 0.92fF
C1839 _330_/A _631_/B 0.44fF
C1840 _607_/X M[12] 0.04fF
C1841 _445_/A _326_/A 1.64fF
C1842 _626_/Y _595_/X 0.03fF
C1843 _573_/A _633_/Y 0.27fF
C1844 _396_/X B[5] 0.01fF
C1845 VPWR _607_/a_493_297# 0.02fF
C1846 _378_/a_664_47# _324_/a_664_47# 0.01fF
C1847 _474_/Y _633_/Y 0.09fF
C1848 _419_/X _383_/X 0.03fF
C1849 _327_/a_493_297# _631_/A 0.01fF
C1850 _461_/a_215_47# _424_/X 0.05fF
C1851 _461_/a_493_297# _423_/X 0.11fF
C1852 _337_/A _475_/A 0.32fF
C1853 _417_/D _512_/a_292_297# 0.02fF
C1854 VPWR _540_/a_250_297# 0.74fF
C1855 _544_/A _565_/a_303_47# 0.03fF
C1856 _627_/D VPWR 8.02fF
C1857 _538_/A _537_/a_77_199# 0.22fF
C1858 VPWR _547_/a_448_47# 0.04fF
C1859 _596_/a_226_47# _626_/Y 0.11fF
C1860 _347_/A _512_/a_292_297# 0.01fF
C1861 _332_/a_68_297# _332_/a_150_297# 0.02fF
C1862 _575_/a_215_47# _547_/X 0.10fF
C1863 _324_/a_558_47# _367_/C 0.24fF
C1864 _583_/X _485_/D 0.03fF
C1865 _601_/Y _607_/a_215_47# 0.24fF
C1866 _606_/Y _607_/a_493_297# 0.08fF
C1867 _612_/Y _610_/Y 0.38fF
C1868 _627_/C _590_/A 0.64fF
C1869 _627_/A _610_/A 0.40fF
C1870 _376_/X _320_/a_161_47# 0.01fF
C1871 _597_/a_215_47# _598_/B 0.29fF
C1872 _632_/a_78_199# _631_/B 0.25fF
C1873 _559_/X _576_/X 2.79fF
C1874 _335_/a_381_47# VPWR 0.34fF
C1875 _432_/B _430_/X 0.01fF
C1876 _602_/Y _504_/X 0.56fF
C1877 _442_/D _530_/X 0.07fF
C1878 _454_/X _511_/X 1.85fF
C1879 _579_/X _530_/X 0.24fF
C1880 _563_/A _380_/A 2.85fF
C1881 input5/a_664_47# _478_/A 0.05fF
C1882 _448_/a_68_297# _447_/B 0.21fF
C1883 _585_/a_109_297# _622_/C 0.02fF
C1884 _567_/B _570_/X 0.07fF
C1885 _477_/a_78_199# _381_/B 0.02fF
C1886 _524_/a_215_47# _489_/X 0.11fF
C1887 _487_/X _547_/X 0.03fF
C1888 _551_/a_226_47# _552_/a_76_199# 0.01fF
C1889 _551_/a_76_199# _552_/a_226_47# 0.01fF
C1890 _322_/A _322_/a_27_47# 0.51fF
C1891 _498_/Y _530_/X 0.01fF
C1892 _513_/a_27_47# _534_/a_80_21# 0.01fF
C1893 _332_/X _366_/a_226_47# 0.30fF
C1894 _486_/B _486_/a_68_297# 0.30fF
C1895 _475_/X _510_/A 0.13fF
C1896 _497_/B _498_/A 0.02fF
C1897 _532_/a_206_369# _557_/B 0.04fF
C1898 _569_/Y _571_/a_584_47# 0.02fF
C1899 _626_/Y _624_/a_76_199# 0.13fF
C1900 _625_/Y _624_/a_489_47# 0.01fF
C1901 _613_/X _616_/A 0.01fF
C1902 _334_/a_27_47# _390_/B 0.31fF
C1903 _379_/a_78_199# VPWR 0.61fF
C1904 _576_/X _616_/B 0.23fF
C1905 _390_/D _537_/a_539_297# 0.03fF
C1906 _490_/X _490_/a_78_199# 0.21fF
C1907 _489_/a_489_413# _489_/a_76_199# 0.12fF
C1908 _424_/X _426_/B 0.01fF
C1909 _625_/a_27_297# _606_/A 0.20fF
C1910 _544_/A _585_/B 0.21fF
C1911 _412_/a_76_199# _458_/a_215_47# 0.01fF
C1912 _567_/B _437_/X 0.40fF
C1913 _520_/a_76_199# VPWR 0.49fF
C1914 _623_/a_489_413# VPWR 0.39fF
C1915 _518_/a_93_21# _381_/B 0.31fF
C1916 _393_/A _631_/Y 1.22fF
C1917 _350_/X _398_/a_489_413# 0.10fF
C1918 _461_/X _462_/a_226_47# 0.53fF
C1919 _616_/Y _606_/A 0.60fF
C1920 _618_/A _625_/a_277_47# 0.06fF
C1921 _436_/A _386_/X 0.04fF
C1922 _613_/X _622_/a_29_53# 0.01fF
C1923 _356_/a_493_297# _452_/A 0.02fF
C1924 B[1] _335_/a_62_47# 0.11fF
C1925 _380_/a_27_47# VPWR 0.59fF
C1926 _349_/a_78_199# _350_/C 0.37fF
C1927 _615_/a_78_199# _573_/Y 0.14fF
C1928 input12/a_381_47# VPWR 0.30fF
C1929 _465_/X _466_/X 1.18fF
C1930 _442_/A _508_/a_227_47# 0.07fF
C1931 _530_/a_76_199# _498_/A 0.02fF
C1932 _390_/D _443_/B 0.03fF
C1933 _579_/a_59_75# VPWR 0.47fF
C1934 _541_/a_78_199# VPWR 0.85fF
C1935 _630_/a_489_413# _629_/X 0.14fF
C1936 _630_/a_76_199# _630_/X 0.22fF
C1937 _479_/a_68_297# VPWR 0.31fF
C1938 _324_/a_62_47# _324_/a_381_47# 0.08fF
C1939 _583_/X A[6] 0.03fF
C1940 _380_/A _351_/a_27_53# 0.16fF
C1941 _616_/B _618_/A 0.02fF
C1942 _426_/B _426_/A 0.60fF
C1943 _422_/a_226_47# _412_/X 0.37fF
C1944 _437_/X _468_/a_78_199# 0.01fF
C1945 _572_/A _609_/a_80_21# 0.11fF
C1946 _549_/X _559_/X 0.46fF
C1947 _550_/X _576_/X 0.01fF
C1948 _387_/a_78_199# _633_/Y 0.12fF
C1949 _487_/X _488_/a_76_199# 0.31fF
C1950 _533_/X _503_/A 0.06fF
C1951 _578_/a_78_199# _533_/X 0.37fF
C1952 _424_/a_76_199# _422_/X 0.38fF
C1953 _424_/a_226_47# _423_/X 0.53fF
C1954 _547_/X _570_/A 0.50fF
C1955 _478_/A _483_/a_93_21# 0.01fF
C1956 _506_/A _479_/B 0.00fF
C1957 _378_/A _324_/a_62_47# 0.12fF
C1958 _473_/a_77_199# _473_/a_323_297# 0.05fF
C1959 _362_/a_489_413# _351_/X 0.07fF
C1960 _460_/X VPWR 1.73fF
C1961 _480_/A _482_/X 0.46fF
C1962 _542_/C _547_/X 0.03fF
C1963 _631_/B _442_/B 0.03fF
C1964 _633_/Y _385_/a_841_47# 0.07fF
C1965 _350_/a_27_297# VPWR 0.43fF
C1966 _332_/X _337_/X 1.98fF
C1967 _608_/a_78_199# _609_/a_80_21# 0.01fF
C1968 _563_/a_27_297# _586_/S 0.20fF
C1969 _485_/A _485_/D 0.04fF
C1970 _587_/A _545_/Y 0.26fF
C1971 _382_/B _382_/a_68_297# 0.30fF
C1972 _570_/a_68_297# _570_/A 0.48fF
C1973 _605_/a_80_21# _602_/Y 0.31fF
C1974 _519_/a_29_53# _519_/X 0.20fF
C1975 _544_/A _447_/X 0.03fF
C1976 _519_/X _417_/D 0.03fF
C1977 _390_/B _337_/A 0.05fF
C1978 _545_/Y _612_/A 0.11fF
C1979 _543_/B _544_/a_381_47# 0.08fF
C1980 _432_/a_68_297# _432_/B 0.33fF
C1981 _436_/A _408_/a_150_297# 0.01fF
C1982 _327_/a_78_199# _445_/A 0.28fF
C1983 _396_/a_256_47# _330_/A 0.04fF
C1984 _386_/X _350_/X 0.05fF
C1985 _455_/X _563_/A 0.03fF
C1986 _609_/a_80_21# _542_/D 0.24fF
C1987 _620_/X _617_/a_113_297# 0.21fF
C1988 _530_/a_76_199# _530_/a_489_413# 0.12fF
C1989 _482_/X _481_/A 1.29fF
C1990 _386_/X _478_/A 0.06fF
C1991 _437_/a_544_297# VPWR 0.01fF
C1992 _633_/A _368_/B 0.12fF
C1993 _455_/X _627_/A 1.41fF
C1994 _563_/D _512_/a_78_199# 0.11fF
C1995 _547_/X _535_/A 0.71fF
C1996 _448_/A _561_/A 0.50fF
C1997 _545_/Y _544_/a_558_47# 0.01fF
C1998 _608_/a_215_47# _572_/A 0.14fF
C1999 _595_/X _593_/A 0.42fF
C2000 _595_/a_227_47# _503_/A 0.03fF
C2001 VPWR _401_/A 0.85fF
C2002 _496_/a_215_47# _460_/X 0.11fF
C2003 _538_/A VPWR 1.54fF
C2004 _510_/X VPWR 1.27fF
C2005 _591_/Y _585_/B 0.18fF
C2006 _482_/a_150_297# _347_/A 0.02fF
C2007 _511_/a_93_21# VPWR 0.43fF
C2008 _567_/B _476_/X 0.03fF
C2009 _627_/A _509_/A 0.03fF
C2010 _326_/a_27_47# _326_/A 0.33fF
C2011 _448_/A B[7] 0.03fF
C2012 _608_/X _503_/A 0.01fF
C2013 _626_/Y _522_/a_226_47# 0.06fF
C2014 A[7] _367_/C 0.03fF
C2015 _551_/X _580_/B 0.01fF
C2016 _630_/a_489_413# _432_/B 0.07fF
C2017 _550_/X _549_/X 1.89fF
C2018 _608_/a_78_199# _608_/a_215_47# 0.26fF
C2019 _443_/a_68_297# VPWR 0.33fF
C2020 _509_/Y _503_/A 0.06fF
C2021 _576_/X _530_/X 0.16fF
C2022 _626_/Y _492_/a_226_47# 0.08fF
C2023 _473_/a_539_297# _472_/Y 0.02fF
C2024 _473_/a_227_47# _471_/Y 0.24fF
C2025 _428_/a_81_21# _428_/a_299_297# 0.21fF
C2026 _356_/a_78_199# _519_/A 0.13fF
C2027 _468_/a_215_47# _503_/A 0.12fF
C2028 _419_/a_76_199# _419_/a_226_47# 0.49fF
C2029 _627_/C _503_/A 0.64fF
C2030 _340_/A _514_/A 0.04fF
C2031 _631_/Y _433_/Y 0.03fF
C2032 _469_/A _485_/D 0.03fF
C2033 _368_/a_68_297# _634_/a_300_297# 0.01fF
C2034 _370_/B _343_/X 0.01fF
C2035 _608_/X _609_/a_209_297# 0.03fF
C2036 _410_/a_27_47# _410_/C 0.18fF
C2037 _594_/X _575_/a_78_199# 0.01fF
C2038 _485_/A A[6] 0.67fF
C2039 _367_/a_27_297# _631_/A 0.32fF
C2040 _532_/a_76_199# _531_/B 0.08fF
C2041 _456_/a_226_47# _456_/X 0.06fF
C2042 _613_/a_77_199# _627_/D 0.48fF
C2043 _464_/A _427_/Y 0.03fF
C2044 _542_/D _627_/a_109_297# 0.01fF
C2045 _573_/A _585_/B 0.61fF
C2046 _487_/a_493_297# _452_/X 0.08fF
C2047 _352_/a_448_47# VPWR 0.03fF
C2048 _385_/a_62_47# _584_/A 0.03fF
C2049 _441_/a_493_297# _454_/X 0.02fF
C2050 _376_/X _542_/D 0.16fF
C2051 _349_/a_78_199# _380_/A 0.17fF
C2052 _634_/a_384_47# _368_/A 0.13fF
C2053 _538_/Y _559_/a_227_297# 0.01fF
C2054 _476_/a_250_297# _471_/Y 0.07fF
C2055 _316_/a_381_47# _316_/a_841_47# 0.03fF
C2056 _316_/a_558_47# _316_/a_664_47# 0.60fF
C2057 _536_/Y _536_/a_109_297# 0.02fF
C2058 _410_/B _346_/A 0.09fF
C2059 _566_/Y _572_/B 0.39fF
C2060 _475_/A VPWR 11.03fF
C2061 _495_/a_76_199# _495_/a_226_47# 0.49fF
C2062 _363_/a_68_297# _363_/a_150_297# 0.02fF
C2063 VPWR _488_/X 1.53fF
C2064 _626_/a_397_297# _626_/Y 0.26fF
C2065 _375_/X _408_/B 0.72fF
C2066 B[1] _510_/A 0.42fF
C2067 _557_/B _558_/a_227_47# 0.18fF
C2068 _530_/a_226_47# _529_/Y 0.55fF
C2069 _410_/B _478_/A 0.07fF
C2070 _611_/a_373_47# _611_/X 0.09fF
C2071 _595_/a_77_199# _595_/a_323_297# 0.05fF
C2072 _436_/A _395_/X 0.12fF
C2073 B[7] _601_/A 0.03fF
C2074 _469_/A _483_/X 0.36fF
C2075 _351_/A _332_/a_68_297# 0.00fF
C2076 _563_/D _631_/B 0.61fF
C2077 _386_/a_62_47# VPWR 0.50fF
C2078 _584_/A _381_/B 0.03fF
C2079 _388_/a_27_47# _411_/A 0.07fF
C2080 B[0] _515_/A 0.03fF
C2081 _561_/A _418_/A 0.10fF
C2082 _491_/a_76_199# VPWR 0.52fF
C2083 _387_/a_215_47# _313_/a_27_47# 0.03fF
C2084 _503_/a_62_47# _627_/A 0.31fF
C2085 _543_/Y _546_/a_226_47# 0.25fF
C2086 _569_/Y _612_/Y 0.03fF
C2087 _593_/Y _598_/A 0.09fF
C2088 _569_/A _627_/A 0.91fF
C2089 _431_/a_556_47# _426_/A 0.02fF
C2090 _633_/a_74_47# VPWR 0.28fF
C2091 _567_/B _402_/a_27_47# 0.32fF
C2092 _371_/B _343_/X 0.04fF
C2093 _597_/a_78_199# VPWR 0.67fF
C2094 _430_/A _430_/X 0.03fF
C2095 _365_/a_299_297# _363_/a_68_297# 0.01fF
C2096 _629_/X _629_/a_68_297# 0.34fF
C2097 _534_/a_80_21# _534_/a_209_297# 0.16fF
C2098 _591_/Y _616_/Y 0.06fF
C2099 _567_/Y _535_/Y 0.17fF
C2100 _626_/Y _521_/X 0.15fF
C2101 _352_/a_448_47# _314_/X 0.22fF
C2102 _311_/a_27_47# _542_/A 0.01fF
C2103 _442_/a_27_47# _631_/Y 0.06fF
C2104 _347_/A _340_/a_27_47# 0.01fF
C2105 _557_/A _557_/Y 0.48fF
C2106 _517_/a_68_297# _517_/X 0.27fF
C2107 _513_/a_27_47# _514_/B 0.20fF
C2108 _603_/a_27_47# _554_/A 0.01fF
C2109 _410_/a_27_47# _445_/X 0.02fF
C2110 _587_/a_27_47# _616_/Y 0.00fF
C2111 _487_/X _480_/A 0.37fF
C2112 _360_/a_226_297# VPWR 0.00fF
C2113 _430_/a_68_297# _432_/B 0.36fF
C2114 _612_/A _617_/a_199_47# 0.01fF
C2115 _542_/A _410_/C 0.31fF
C2116 _610_/A _621_/a_215_47# 0.10fF
C2117 _549_/X _530_/X 0.17fF
C2118 _471_/Y _509_/Y 0.02fF
C2119 _455_/a_222_93# _419_/X 0.01fF
C2120 M[0] _552_/a_76_199# 0.05fF
C2121 _557_/A _467_/Y 0.43fF
C2122 M[7] VPWR 1.00fF
C2123 _413_/X _419_/a_226_297# 0.02fF
C2124 _494_/a_226_47# VPWR 0.08fF
C2125 _556_/Y _558_/a_227_47# 0.10fF
C2126 _455_/a_79_199# _455_/X 0.29fF
C2127 _455_/a_222_93# _413_/X 0.03fF
C2128 _411_/B _410_/C 0.07fF
C2129 _469_/A A[6] 0.01fF
C2130 _469_/a_62_47# _584_/A 0.07fF
C2131 _510_/A _383_/X 0.03fF
C2132 M[6] _621_/X 0.83fF
C2133 _365_/a_81_21# _365_/a_299_297# 0.21fF
C2134 _386_/A _385_/a_62_47# 0.31fF
C2135 _491_/a_226_47# _490_/X 0.53fF
C2136 _627_/A _627_/D 1.28fF
C2137 _485_/a_27_47# _542_/D 0.36fF
C2138 _395_/X _350_/X 0.21fF
C2139 _563_/a_27_297# _563_/a_109_297# 0.02fF
C2140 _352_/X _361_/X 0.78fF
C2141 _627_/C _627_/a_205_297# 0.01fF
C2142 _553_/a_78_199# _525_/X 0.40fF
C2143 _627_/C _590_/a_150_297# 0.01fF
C2144 VPWR _617_/a_113_297# 0.57fF
C2145 _448_/A VPWR 1.76fF
C2146 _483_/X _489_/a_76_199# 0.21fF
C2147 _587_/A _458_/X 0.05fF
C2148 B[1] _631_/A 0.42fF
C2149 M[9] _542_/D 0.10fF
C2150 _508_/a_227_47# _509_/A 0.04fF
C2151 _495_/a_76_199# _494_/X 0.34fF
C2152 _495_/a_226_47# _468_/X 0.31fF
C2153 _487_/X _481_/A 0.36fF
C2154 _417_/D _480_/Y 0.06fF
C2155 _426_/A _629_/B 0.38fF
C2156 _595_/a_539_297# _570_/X 0.02fF
C2157 _595_/a_227_47# _566_/Y 0.07fF
C2158 _386_/A _381_/B 1.13fF
C2159 _412_/X _437_/a_79_199# 0.01fF
C2160 _635_/Y _370_/B 0.13fF
C2161 _412_/a_489_413# _408_/X 0.17fF
C2162 _482_/a_68_297# _563_/D 0.30fF
C2163 _534_/a_209_297# _530_/X 0.14fF
C2164 _487_/X _633_/Y 0.07fF
C2165 _359_/a_68_297# _381_/B 0.01fF
C2166 _411_/a_68_297# _411_/a_150_297# 0.02fF
C2167 _406_/A _420_/X 2.10fF
C2168 _349_/a_292_297# _419_/X 0.02fF
C2169 _573_/A _572_/B 0.17fF
C2170 _543_/B _469_/a_841_47# 0.01fF
C2171 _431_/a_76_199# _431_/a_226_47# 0.49fF
C2172 VPWR _511_/X 2.75fF
C2173 _431_/a_489_413# _478_/A 0.09fF
C2174 _516_/A _417_/D 0.10fF
C2175 _439_/X _567_/B 0.16fF
C2176 _578_/a_493_297# VPWR 0.01fF
C2177 _519_/A _486_/A 0.01fF
C2178 _443_/B _631_/Y 0.25fF
C2179 _623_/a_226_47# M[6] 0.07fF
C2180 A[6] _489_/a_76_199# 0.01fF
C2181 _417_/D _539_/A 0.29fF
C2182 _631_/Y _316_/a_664_47# 0.08fF
C2183 _381_/C _481_/A 2.26fF
C2184 _473_/a_77_199# VPWR 0.92fF
C2185 _626_/Y _575_/X 0.09fF
C2186 _411_/B _445_/X 0.03fF
C2187 _584_/A _542_/A 0.15fF
C2188 output21/a_27_47# _626_/a_397_297# 0.03fF
C2189 _583_/X _581_/B 0.61fF
C2190 _432_/A VPWR 1.25fF
C2191 _347_/A _539_/A 0.66fF
C2192 _516_/A _347_/A 0.55fF
C2193 _390_/B VPWR 11.47fF
C2194 _520_/X _469_/X 0.19fF
C2195 _542_/C _480_/A 0.29fF
C2196 VPWR _601_/A 2.14fF
C2197 _557_/A _606_/A 0.35fF
C2198 _613_/a_323_297# _590_/A 0.04fF
C2199 _455_/a_79_199# _452_/A 0.18fF
C2200 _350_/a_277_297# _350_/C 0.01fF
C2201 _383_/X _631_/A 0.67fF
C2202 _416_/a_215_47# _561_/A 0.03fF
C2203 _513_/A _417_/a_197_47# 0.03fF
C2204 _599_/A _598_/B 0.01fF
C2205 _493_/X VPWR 2.96fF
C2206 _403_/a_27_47# _486_/X 0.10fF
C2207 _635_/Y _371_/B 0.19fF
C2208 _445_/A _326_/a_27_47# 0.29fF
C2209 _625_/Y _624_/X 0.51fF
C2210 _439_/X _468_/a_78_199# 0.28fF
C2211 _417_/a_109_47# _542_/A 0.02fF
C2212 _504_/a_227_47# _471_/Y 0.07fF
C2213 _519_/X _547_/a_79_199# 0.23fF
C2214 _370_/A _635_/a_27_413# 0.09fF
C2215 _628_/a_382_297# _625_/Y 0.05fF
C2216 _418_/A VPWR 0.63fF
C2217 _587_/A _622_/C 0.02fF
C2218 _375_/a_79_199# _481_/A 0.01fF
C2219 _519_/A _332_/a_68_297# 0.30fF
C2220 _606_/Y _601_/A 0.04fF
C2221 M[0] output17/a_27_47# 0.61fF
C2222 _588_/A _593_/Y 0.01fF
C2223 _419_/X _458_/a_78_199# 0.01fF
C2224 _468_/X _494_/X 1.52fF
C2225 _350_/a_27_297# _563_/A 0.44fF
C2226 _612_/A _622_/C 0.91fF
C2227 _467_/Y _527_/Y 0.24fF
C2228 _474_/Y _476_/a_250_297# 0.06fF
C2229 _542_/C _481_/A 0.34fF
C2230 _549_/a_489_413# VPWR 0.39fF
C2231 _374_/X _399_/a_78_199# 0.02fF
C2232 _456_/a_556_47# VPWR 0.00fF
C2233 _420_/X _350_/C 0.04fF
C2234 _424_/a_226_297# VPWR 0.00fF
C2235 _453_/a_256_47# _542_/D 0.04fF
C2236 _525_/a_226_297# _523_/X 0.01fF
C2237 output19/a_27_47# VPWR 0.66fF
C2238 input3/a_62_47# _485_/D 0.05fF
C2239 _469_/A _549_/a_226_47# 0.00fF
C2240 _465_/X _467_/a_397_297# 0.12fF
C2241 _386_/X _381_/B 0.56fF
C2242 _408_/B _337_/B 0.01fF
C2243 _591_/Y _627_/C 0.23fF
C2244 _595_/a_77_199# VPWR 0.89fF
C2245 _580_/a_68_297# _581_/B 0.27fF
C2246 _567_/Y A[3] 0.03fF
C2247 _519_/A _328_/A 0.69fF
C2248 _612_/A _618_/Y 0.45fF
C2249 _390_/B _501_/Y 0.60fF
C2250 _542_/B _478_/a_197_47# 0.08fF
C2251 _629_/A _630_/a_76_199# 0.06fF
C2252 _328_/B VPWR 1.11fF
C2253 _340_/A _512_/a_215_47# 0.16fF
C2254 _625_/Y _622_/C 0.05fF
C2255 B[0] A[3] 0.05fF
C2256 _623_/X _627_/B 0.41fF
C2257 _602_/Y _556_/A 0.08fF
C2258 _420_/X _367_/C 0.12fF
C2259 _386_/A _542_/A 0.02fF
C2260 M[5] _374_/X 0.06fF
C2261 _504_/a_227_47# _504_/X 0.04fF
C2262 _471_/A VPWR 1.70fF
C2263 _476_/X _476_/a_93_21# 0.13fF
C2264 _411_/A _350_/C 0.02fF
C2265 _411_/B _386_/A 0.03fF
C2266 _545_/Y _433_/Y 0.02fF
C2267 _586_/S _545_/Y 0.05fF
C2268 _568_/a_539_297# _546_/X 0.04fF
C2269 _506_/A _478_/A 0.56fF
C2270 input8/a_27_47# A[7] 0.40fF
C2271 _623_/X _620_/X 0.36fF
C2272 _611_/a_109_297# _591_/Y 0.05fF
C2273 _533_/a_77_199# _503_/A 0.50fF
C2274 _511_/a_250_297# _433_/Y 0.02fF
C2275 _424_/a_76_199# _406_/Y 0.02fF
C2276 _459_/a_226_47# _457_/X 0.35fF
C2277 _538_/A _627_/A 0.26fF
C2278 _601_/Y _618_/Y 0.19fF
C2279 _448_/B _453_/a_250_297# 0.01fF
C2280 _510_/X _627_/A 0.18fF
C2281 _474_/Y _468_/a_215_47# 0.01fF
C2282 _390_/D _538_/Y 1.14fF
C2283 _510_/A _438_/a_150_297# 0.01fF
C2284 _633_/Y _419_/X 0.03fF
C2285 _375_/X _337_/B 0.13fF
C2286 _424_/X _406_/A 0.02fF
C2287 _432_/B _398_/X 0.01fF
C2288 _461_/a_215_47# _407_/Y 0.12fF
C2289 _469_/A input16/a_27_47# 0.22fF
C2290 _446_/X _472_/B 0.05fF
C2291 _543_/A _610_/A 0.01fF
C2292 _623_/X B[7] 1.48fF
C2293 _417_/D _340_/A 0.43fF
C2294 _585_/B _539_/X 0.23fF
C2295 _417_/D _479_/A 0.12fF
C2296 _604_/a_80_21# _604_/a_209_47# 0.04fF
C2297 B[2] _606_/A 0.03fF
C2298 _632_/a_78_199# _320_/a_161_47# 0.02fF
C2299 _619_/a_109_297# VPWR 0.01fF
C2300 _504_/a_77_199# _504_/a_323_297# 0.05fF
C2301 _426_/A _399_/a_78_199# 0.21fF
C2302 VPWR _524_/X 1.39fF
C2303 _467_/Y _531_/A 0.41fF
C2304 _347_/A _479_/A 0.01fF
C2305 _621_/a_78_199# _621_/a_215_47# 0.26fF
C2306 _531_/a_109_297# _558_/X 0.08fF
C2307 _376_/X _383_/a_76_199# 0.42fF
C2308 _347_/A _340_/A 2.48fF
C2309 _369_/a_226_47# B[5] 0.06fF
C2310 _371_/B _370_/B 0.13fF
C2311 _534_/a_209_297# _514_/B 0.03fF
C2312 _623_/X _589_/a_226_47# 0.06fF
C2313 _370_/a_68_297# B[5] 0.11fF
C2314 _563_/A _475_/A 0.26fF
C2315 _487_/X _521_/a_78_199# 0.13fF
C2316 _415_/a_27_47# _542_/A 0.10fF
C2317 _469_/A _570_/X 0.63fF
C2318 _554_/B _554_/a_68_297# 0.32fF
C2319 _606_/Y _619_/a_109_297# 0.07fF
C2320 _330_/A _352_/X 0.06fF
C2321 _416_/a_215_47# VPWR 0.04fF
C2322 _455_/X _490_/a_493_297# 0.09fF
C2323 _486_/A _486_/X 0.03fF
C2324 _397_/a_226_47# _397_/a_489_413# 0.02fF
C2325 _397_/a_76_199# _397_/a_226_297# 0.01fF
C2326 _436_/A _412_/a_489_413# 0.11fF
C2327 _459_/a_226_47# _459_/X 0.05fF
C2328 _437_/a_79_199# _411_/X 0.31fF
C2329 _445_/A _387_/a_215_47# 0.05fF
C2330 _573_/Y _574_/a_81_21# 0.39fF
C2331 _447_/X _519_/C 0.27fF
C2332 _485_/D _547_/X 2.00fF
C2333 _426_/A M[5] 0.08fF
C2334 _596_/a_76_199# _594_/X 0.43fF
C2335 _430_/A _430_/a_68_297# 0.30fF
C2336 _513_/A _486_/A 0.05fF
C2337 _627_/A _475_/A 0.12fF
C2338 _386_/X _542_/A 0.28fF
C2339 _604_/X _530_/X 0.06fF
C2340 _390_/D _486_/X 0.03fF
C2341 _475_/A _438_/a_68_297# 0.29fF
C2342 _542_/B _479_/B 0.02fF
C2343 _410_/a_27_47# _410_/B 0.39fF
C2344 _407_/Y _426_/B 0.03fF
C2345 _342_/X _328_/B 0.26fF
C2346 _423_/a_78_199# _423_/a_215_47# 0.26fF
C2347 _417_/D _521_/a_493_297# 0.02fF
C2348 _488_/a_226_47# _520_/X 0.23fF
C2349 _355_/a_161_47# _442_/A 0.03fF
C2350 _411_/B _386_/X 0.61fF
C2351 VPWR _604_/a_80_21# 0.32fF
C2352 _426_/A _428_/X 0.41fF
C2353 _380_/A _363_/A 0.03fF
C2354 _485_/D _570_/a_68_297# 0.05fF
C2355 _504_/a_77_199# VPWR 0.89fF
C2356 _380_/A _420_/X 0.03fF
C2357 _441_/a_493_297# VPWR 0.01fF
C2358 _562_/a_493_297# _584_/A 0.01fF
C2359 _477_/a_78_199# _539_/A 0.17fF
C2360 _493_/a_78_199# _493_/a_215_47# 0.26fF
C2361 _516_/A _477_/a_78_199# 0.31fF
C2362 _586_/a_535_374# _433_/Y 0.00fF
C2363 _515_/Y _570_/A 0.51fF
C2364 _503_/a_381_47# _503_/a_558_47# 0.32fF
C2365 _350_/C _409_/a_78_199# 0.40fF
C2366 _371_/A _373_/Y 0.21fF
C2367 _508_/a_323_297# _507_/Y 0.01fF
C2368 _474_/Y _504_/a_227_47# 0.05fF
C2369 _563_/B _519_/C 0.75fF
C2370 _603_/a_27_47# _579_/X 0.08fF
C2371 _420_/X _421_/a_489_413# 0.14fF
C2372 _570_/X _559_/a_227_47# 0.03fF
C2373 _626_/Y M[14] 0.18fF
C2374 _586_/S _586_/a_535_374# 0.02fF
C2375 _436_/A _391_/A 0.03fF
C2376 _503_/A _469_/X 0.94fF
C2377 _534_/a_209_47# _381_/B 0.01fF
C2378 _543_/Y _542_/C 0.43fF
C2379 _542_/C _515_/Y 0.05fF
C2380 _487_/X _585_/B 0.16fF
C2381 _538_/A _537_/a_227_47# 0.04fF
C2382 _544_/A _417_/A 0.30fF
C2383 VPWR _439_/a_226_47# 0.11fF
C2384 _542_/B B[0] 0.05fF
C2385 _390_/D _454_/X 0.03fF
C2386 _464_/A _467_/Y 0.01fF
C2387 M[14] _467_/a_109_47# 0.01fF
C2388 _371_/A VPWR 0.99fF
C2389 _469_/A _590_/B 0.01fF
C2390 input3/a_381_47# _606_/A 0.18fF
C2391 _595_/X _598_/A 0.01fF
C2392 _453_/a_93_21# _453_/a_250_297# 0.50fF
C2393 _616_/B _593_/Y 0.26fF
C2394 _625_/Y _612_/A 2.11fF
C2395 _378_/A _447_/B 0.27fF
C2396 _420_/a_79_199# _420_/a_222_93# 0.51fF
C2397 _609_/a_209_297# _469_/X 0.07fF
C2398 _413_/X _413_/a_68_297# 0.27fF
C2399 _605_/a_80_21# _557_/A 0.31fF
C2400 _447_/a_68_297# _542_/D 0.20fF
C2401 VPWR _361_/a_226_47# 0.06fF
C2402 input3/a_841_47# _616_/B 0.01fF
C2403 _573_/Y VPWR 1.67fF
C2404 _515_/Y _535_/A 0.46fF
C2405 _596_/a_226_47# _598_/A 0.05fF
C2406 _544_/a_381_47# VPWR 0.30fF
C2407 _623_/X VPWR 4.47fF
C2408 _384_/X VPWR 2.52fF
C2409 _314_/a_68_297# _314_/a_150_297# 0.02fF
C2410 _411_/B _410_/B 1.06fF
C2411 M[2] _368_/B 0.18fF
C2412 _544_/a_381_47# _544_/a_664_47# 0.09fF
C2413 _572_/A A[3] 0.03fF
C2414 _458_/X _433_/Y 0.03fF
C2415 _604_/X _557_/B 0.15fF
C2416 _391_/A _350_/X 0.71fF
C2417 _579_/X _554_/A 0.00fF
C2418 _335_/a_62_47# _633_/Y 0.10fF
C2419 _431_/a_76_199# _431_/X 0.24fF
C2420 _478_/A _432_/X 0.03fF
C2421 M[13] _583_/X 0.08fF
C2422 _487_/X _447_/X 0.01fF
C2423 _567_/B _455_/X 0.50fF
C2424 _523_/a_226_47# _521_/X 0.01fF
C2425 _585_/B _570_/A 0.24fF
C2426 _563_/A _390_/B 0.12fF
C2427 _379_/a_215_47# _452_/A 0.03fF
C2428 _627_/A _511_/X 0.03fF
C2429 _337_/a_68_297# _337_/A 0.32fF
C2430 _380_/A _374_/X 0.19fF
C2431 _436_/A _330_/A 0.23fF
C2432 _382_/B _542_/D 0.96fF
C2433 _585_/B _508_/a_77_199# 0.34fF
C2434 _491_/X VPWR 1.05fF
C2435 _531_/B _530_/X 0.26fF
C2436 _496_/a_292_297# VPWR 0.01fF
C2437 _480_/Y _410_/C 0.75fF
C2438 _444_/Y VPWR 1.85fF
C2439 _554_/X _582_/a_109_297# 0.01fF
C2440 _627_/A _473_/a_77_199# 0.06fF
C2441 _490_/a_78_199# _490_/a_292_297# 0.03fF
C2442 _471_/Y _469_/X 0.72fF
C2443 _352_/X _442_/B 0.01fF
C2444 _404_/a_558_47# _503_/A 0.11fF
C2445 VPWR _559_/a_227_297# 0.01fF
C2446 _457_/a_76_199# _457_/a_226_47# 0.49fF
C2447 _549_/X _551_/a_226_297# 0.01fF
C2448 _627_/A _390_/B 0.08fF
C2449 _368_/B _332_/X 0.23fF
C2450 _628_/a_382_297# _433_/Y 0.14fF
C2451 _610_/Y _617_/a_199_47# 0.01fF
C2452 input10/a_27_47# VPWR 0.54fF
C2453 _487_/X _563_/B 0.29fF
C2454 _381_/C _447_/X 0.12fF
C2455 _627_/A _609_/a_303_47# 0.01fF
C2456 _386_/a_841_47# _570_/A 0.07fF
C2457 _433_/a_109_297# _431_/X 0.01fF
C2458 _433_/a_109_47# _432_/X 0.74fF
C2459 _464_/A _427_/A 1.06fF
C2460 _375_/a_79_199# _359_/X 0.35fF
C2461 _503_/A _546_/X 0.03fF
C2462 _567_/Y _548_/a_556_47# 0.05fF
C2463 _574_/X _546_/X 0.35fF
C2464 _335_/a_381_47# _335_/a_841_47# 0.03fF
C2465 _335_/a_558_47# _335_/a_664_47# 0.60fF
C2466 _448_/B _449_/A 0.01fF
C2467 _631_/B _503_/A 0.12fF
C2468 _477_/a_78_199# _479_/A 0.21fF
C2469 _556_/Y _604_/X 0.74fF
C2470 _340_/A _477_/a_78_199# 0.25fF
C2471 _329_/a_76_199# VPWR 0.48fF
C2472 _539_/A _410_/C 0.41fF
C2473 _585_/B _535_/A 0.78fF
C2474 VPWR _394_/a_841_47# 0.40fF
C2475 B[0] _563_/D 0.16fF
C2476 _503_/A _570_/a_150_297# 0.02fF
C2477 _410_/B _470_/a_303_47# 0.07fF
C2478 _360_/X _332_/X 0.16fF
C2479 _627_/C _519_/C 0.98fF
C2480 _417_/D _418_/a_150_297# 0.02fF
C2481 _519_/a_183_297# _563_/B 0.03fF
C2482 _400_/a_303_47# _391_/B 0.01fF
C2483 _381_/C _563_/B 1.92fF
C2484 _390_/D _549_/a_556_47# 0.02fF
C2485 _433_/Y _622_/C 0.16fF
C2486 _562_/a_78_199# _451_/a_27_47# 0.00fF
C2487 _349_/a_78_199# _475_/A 0.28fF
C2488 _528_/a_299_297# VPWR 0.68fF
C2489 _553_/a_215_47# _554_/B 0.13fF
C2490 _330_/A _350_/X 0.03fF
C2491 _479_/A _518_/a_93_21# 0.01fF
C2492 _526_/a_76_199# _526_/a_226_47# 0.49fF
C2493 _485_/A _317_/a_27_47# 0.22fF
C2494 _559_/a_77_199# _559_/a_227_47# 0.24fF
C2495 _563_/D _408_/X 0.05fF
C2496 _454_/X _316_/a_558_47# 0.08fF
C2497 _328_/A _337_/A 0.02fF
C2498 _627_/A _595_/a_77_199# 0.65fF
C2499 _586_/S _622_/C 0.57fF
C2500 _566_/Y _469_/X 0.86fF
C2501 _361_/a_489_413# _361_/a_76_199# 0.12fF
C2502 _390_/D _537_/a_77_199# 0.19fF
C2503 _335_/a_558_47# _519_/A 0.29fF
C2504 _471_/A _470_/a_80_21# 0.20fF
C2505 _387_/a_493_297# VPWR 0.01fF
C2506 _595_/X _588_/A 0.38fF
C2507 _549_/a_226_297# _540_/X 0.02fF
C2508 _549_/a_489_413# _548_/X 0.14fF
C2509 _342_/a_68_297# _342_/a_150_297# 0.02fF
C2510 _569_/A _567_/B 0.08fF
C2511 _329_/a_76_199# _314_/X 0.45fF
C2512 _485_/a_27_47# _542_/A 0.23fF
C2513 _356_/a_78_199# VPWR 0.65fF
C2514 _531_/B _557_/B 0.24fF
C2515 _627_/A _471_/A 0.63fF
C2516 _561_/A _486_/A 0.47fF
C2517 _596_/a_489_413# _599_/Y 0.00fF
C2518 _514_/B _514_/A 0.83fF
C2519 _440_/a_489_413# VPWR 0.39fF
C2520 _403_/a_27_47# VPWR 0.72fF
C2521 _379_/a_78_199# _379_/a_215_47# 0.26fF
C2522 _420_/X _452_/A 0.09fF
C2523 _515_/Y _518_/a_256_47# 0.02fF
C2524 _570_/B _535_/Y 0.06fF
C2525 VPWR _399_/a_292_297# 0.01fF
C2526 _569_/Y _545_/Y 0.03fF
C2527 _530_/X _554_/B 0.13fF
C2528 _591_/A _599_/Y 0.88fF
C2529 _385_/a_62_47# _394_/a_381_47# 0.01fF
C2530 _408_/B _408_/a_68_297# 0.30fF
C2531 _516_/A _584_/A 0.90fF
C2532 _418_/X _324_/a_381_47# 0.18fF
C2533 _418_/A _324_/a_558_47# 0.01fF
C2534 _390_/D B[7] 0.03fF
C2535 _612_/Y B[7] 0.18fF
C2536 _329_/a_76_199# _329_/a_489_413# 0.12fF
C2537 VPWR A[0] 0.55fF
C2538 _544_/A _546_/X 0.06fF
C2539 _510_/A _481_/A 0.15fF
C2540 _520_/a_76_199# _520_/a_226_297# 0.01fF
C2541 _520_/a_226_47# _520_/a_489_413# 0.02fF
C2542 _383_/a_76_199# _383_/a_226_297# 0.01fF
C2543 _383_/a_226_47# _383_/a_489_413# 0.02fF
C2544 _571_/a_250_297# _381_/B 0.04fF
C2545 _420_/X _421_/X 0.21fF
C2546 _610_/Y _622_/C 0.04fF
C2547 _406_/B VPWR 1.33fF
C2548 _487_/X _537_/a_323_297# 0.02fF
C2549 _417_/A B[5] 0.50fF
C2550 _462_/X _461_/X 0.17fF
C2551 _378_/A _418_/X 0.28fF
C2552 _563_/a_27_297# _451_/A 0.02fF
C2553 _510_/A _633_/Y 2.52fF
C2554 _529_/a_109_297# VPWR 0.01fF
C2555 _599_/Y _624_/a_206_369# 0.06fF
C2556 _436_/A _442_/B 0.45fF
C2557 _612_/Y _589_/a_226_47# 0.07fF
C2558 _449_/A _453_/a_93_21# 0.47fF
C2559 _460_/a_226_47# _460_/X 0.05fF
C2560 _352_/a_79_199# _328_/a_68_297# 0.01fF
C2561 _381_/B _515_/A 1.08fF
C2562 _386_/A _480_/Y 0.22fF
C2563 _557_/A _531_/a_109_297# 0.03fF
C2564 _523_/X _511_/X 0.06fF
C2565 _500_/a_78_199# _500_/a_215_47# 0.26fF
C2566 _574_/X _548_/a_76_199# 0.00fF
C2567 _485_/A _367_/C 0.00fF
C2568 _533_/X _552_/a_226_47# 0.33fF
C2569 _551_/X _552_/a_76_199# 0.22fF
C2570 _633_/Y _485_/D 0.03fF
C2571 _487_/X _627_/C 0.52fF
C2572 _396_/X _631_/A 0.23fF
C2573 _542_/B _542_/D 0.10fF
C2574 _396_/a_346_47# _386_/X 0.06fF
C2575 _631_/B _391_/B 0.51fF
C2576 output22/a_27_47# _466_/X 0.01fF
C2577 _419_/a_226_47# _418_/X 0.53fF
C2578 _385_/a_381_47# _385_/a_558_47# 0.32fF
C2579 input12/a_381_47# input12/a_841_47# 0.03fF
C2580 input12/a_558_47# input12/a_664_47# 0.60fF
C2581 VPWR _469_/a_841_47# 0.34fF
C2582 _568_/a_77_199# _568_/a_323_297# 0.05fF
C2583 _340_/A _410_/C 0.01fF
C2584 _455_/a_222_93# _418_/B 0.25fF
C2585 VPWR _555_/a_215_297# 0.37fF
C2586 _454_/X _628_/Y 0.47fF
C2587 _417_/D _448_/B 0.70fF
C2588 _396_/a_250_297# _391_/a_68_297# 0.03fF
C2589 _375_/X _359_/B 0.13fF
C2590 _485_/A _442_/A 1.67fF
C2591 _623_/X _613_/a_77_199# 0.15fF
C2592 _566_/Y _546_/X 0.60fF
C2593 _570_/X _547_/X 0.25fF
C2594 _381_/B _535_/Y 0.05fF
C2595 _498_/A _530_/X 0.01fF
C2596 _474_/Y _469_/X 0.40fF
C2597 _541_/a_78_199# _541_/a_215_47# 0.26fF
C2598 B[4] _374_/X 0.06fF
C2599 _516_/A _386_/A 0.61fF
C2600 _386_/A _539_/A 0.17fF
C2601 _454_/X _631_/Y 5.24fF
C2602 _481_/a_27_47# _486_/X 0.10fF
C2603 _468_/a_215_47# _438_/X 0.12fF
C2604 _417_/D _530_/X 0.05fF
C2605 _504_/a_77_199# _627_/A 0.45fF
C2606 M[0] _606_/A 0.05fF
C2607 _381_/C _627_/C 0.47fF
C2608 _412_/a_76_199# _412_/a_226_47# 0.49fF
C2609 _570_/X _570_/a_68_297# 0.27fF
C2610 _480_/Y _483_/a_93_21# 0.32fF
C2611 _633_/Y _483_/X 0.35fF
C2612 _367_/a_27_297# _367_/C 0.55fF
C2613 _631_/A _481_/A 0.48fF
C2614 _532_/a_206_369# _498_/Y 0.06fF
C2615 _442_/B _350_/X 0.22fF
C2616 _347_/A _530_/X 0.05fF
C2617 _480_/A A[6] 0.04fF
C2618 _451_/A _628_/Y 0.24fF
C2619 _633_/Y _631_/A 0.44fF
C2620 _587_/A _433_/Y 0.78fF
C2621 _544_/A _482_/a_68_297# 0.00fF
C2622 _543_/A _541_/a_78_199# 0.21fF
C2623 _433_/Y _439_/a_489_413# 0.02fF
C2624 _442_/B _346_/A 0.43fF
C2625 _454_/X _452_/X 0.04fF
C2626 _360_/X input13/a_27_47# 0.01fF
C2627 _540_/a_256_47# _486_/X 0.01fF
C2628 _542_/B _478_/A 0.31fF
C2629 _487_/a_292_297# VPWR 0.01fF
C2630 _442_/B _478_/A 0.35fF
C2631 _422_/a_226_47# _422_/X 0.05fF
C2632 _586_/S _612_/A 0.09fF
C2633 _337_/a_68_297# VPWR 0.29fF
C2634 _442_/B _369_/a_489_413# 0.09fF
C2635 _381_/a_27_47# _381_/B 0.37fF
C2636 _376_/X _420_/a_222_93# 0.03fF
C2637 VPWR _486_/A 0.75fF
C2638 _567_/B _460_/X 0.06fF
C2639 _350_/a_27_297# _350_/a_277_297# 0.05fF
C2640 A[6] _481_/A 0.05fF
C2641 _527_/B _602_/Y 0.00fF
C2642 _563_/a_27_297# _627_/B 0.02fF
C2643 _549_/X _554_/A 0.01fF
C2644 _543_/a_109_297# _543_/Y 0.03fF
C2645 _340_/A _584_/A 1.21fF
C2646 _463_/a_489_413# _626_/Y 0.09fF
C2647 _612_/Y VPWR 2.42fF
C2648 _386_/X _480_/Y 0.29fF
C2649 _568_/a_323_297# _566_/A 0.01fF
C2650 _491_/a_489_413# _490_/a_78_199# 0.01fF
C2651 _557_/A _556_/A 0.02fF
C2652 _390_/D VPWR 7.30fF
C2653 _510_/a_68_297# _510_/A 0.35fF
C2654 _568_/a_539_297# _567_/Y 0.03fF
C2655 _633_/Y A[6] 0.11fF
C2656 _625_/Y _433_/Y 0.43fF
C2657 _570_/B A[3] 0.16fF
C2658 _475_/a_68_297# _475_/A 0.35fF
C2659 _571_/a_256_47# _469_/X 0.02fF
C2660 _625_/Y _586_/S 0.20fF
C2661 _623_/X _627_/A 0.16fF
C2662 _616_/a_109_297# _616_/A 0.02fF
C2663 _513_/A _355_/A 0.60fF
C2664 _436_/A _563_/D 0.17fF
C2665 _362_/a_76_199# _371_/B 0.18fF
C2666 _519_/A _447_/B 2.27fF
C2667 _536_/a_109_297# _530_/X 0.02fF
C2668 _519_/X _485_/a_27_47# 0.02fF
C2669 _542_/A _515_/A 0.59fF
C2670 _551_/X output17/a_27_47# 0.02fF
C2671 B[1] _350_/C 0.10fF
C2672 M[3] B[5] 0.40fF
C2673 _584_/A _588_/A 0.36fF
C2674 _543_/B _565_/a_80_21# 0.68fF
C2675 _380_/A _485_/A 0.98fF
C2676 _404_/a_62_47# _544_/a_381_47# 0.02fF
C2677 _410_/B _340_/a_27_47# 0.10fF
C2678 _595_/X _616_/B 0.01fF
C2679 _628_/a_734_297# _628_/Y 0.33fF
C2680 _466_/a_215_47# _430_/X 0.13fF
C2681 _543_/B _545_/Y 0.19fF
C2682 _382_/B _383_/a_76_199# 0.01fF
C2683 _635_/Y _635_/a_384_47# 0.01fF
C2684 _406_/A _405_/a_109_297# 0.01fF
C2685 VPWR _332_/a_68_297# 0.34fF
C2686 _563_/D _542_/D 0.06fF
C2687 _563_/a_27_297# _561_/A 0.01fF
C2688 _595_/X _571_/a_93_21# 0.03fF
C2689 B[0] _520_/X 0.55fF
C2690 _490_/a_78_199# _454_/X 0.01fF
C2691 _632_/a_215_47# VPWR 0.07fF
C2692 _573_/Y _548_/X 0.02fF
C2693 _386_/X _539_/A 0.27fF
C2694 _516_/A _386_/X 1.85fF
C2695 _504_/a_227_47# _438_/X 0.00fF
C2696 _362_/a_226_47# _361_/a_226_47# 0.02fF
C2697 _533_/a_227_47# _503_/A 0.19fF
C2698 _519_/A _376_/a_68_297# 0.14fF
C2699 _463_/a_226_47# _462_/X 0.54fF
C2700 _463_/a_489_413# _406_/Y 0.16fF
C2701 input2/a_27_47# VPWR 0.71fF
C2702 _610_/Y _612_/A 2.63fF
C2703 _355_/A _454_/X 0.09fF
C2704 _444_/Y _470_/a_80_21# 0.41fF
C2705 _600_/a_27_297# _601_/A 0.25fF
C2706 _567_/B _538_/A 0.01fF
C2707 _596_/a_226_47# _616_/B 0.06fF
C2708 _567_/B _401_/A 0.57fF
C2709 _565_/a_80_21# _565_/a_209_297# 0.16fF
C2710 _500_/a_78_199# _500_/a_292_297# 0.03fF
C2711 _359_/A _383_/X 0.06fF
C2712 _629_/X _629_/B 0.14fF
C2713 input5/a_381_47# input5/a_664_47# 0.09fF
C2714 _444_/Y _627_/A 0.01fF
C2715 B[1] _367_/C 0.02fF
C2716 _356_/a_215_47# _359_/A 0.01fF
C2717 _436_/X _436_/a_68_297# 0.27fF
C2718 _577_/a_226_47# _559_/X 0.23fF
C2719 _577_/a_76_199# _576_/X 0.22fF
C2720 _328_/A VPWR 1.77fF
C2721 _523_/X _524_/X 2.64fF
C2722 _390_/D _559_/a_539_297# 0.03fF
C2723 _627_/A _559_/a_227_297# 0.04fF
C2724 _420_/a_448_47# _320_/a_161_47# 0.03fF
C2725 _406_/A _407_/Y 0.01fF
C2726 output27/a_27_47# _629_/B 0.30fF
C2727 _382_/B _381_/B 0.02fF
C2728 _437_/a_79_199# _408_/X 0.01fF
C2729 _628_/Y _627_/B 0.47fF
C2730 VPWR _324_/a_62_47# 0.48fF
C2731 _469_/a_381_47# _469_/a_558_47# 0.32fF
C2732 _386_/A _340_/A 0.03fF
C2733 M[8] A[1] 0.04fF
C2734 _469_/A _610_/A 0.68fF
C2735 _515_/Y _485_/D 0.99fF
C2736 _479_/a_150_297# _486_/X 0.01fF
C2737 _386_/A _479_/A 0.22fF
C2738 _625_/Y _610_/Y 0.13fF
C2739 _587_/A _537_/a_539_297# 0.04fF
C2740 _351_/A _350_/B 0.43fF
C2741 _383_/X _350_/C 0.90fF
C2742 _386_/a_664_47# _479_/a_68_297# 0.01fF
C2743 A[3] _381_/B 0.17fF
C2744 _568_/a_227_47# _585_/B 0.03fF
C2745 _563_/D _346_/A 0.33fF
C2746 _465_/a_27_297# _464_/A 0.36fF
C2747 _542_/a_27_47# _514_/a_68_297# 0.01fF
C2748 _616_/A _624_/a_206_369# 0.10fF
C2749 _616_/B _624_/a_76_199# 0.12fF
C2750 _616_/Y _624_/a_585_369# 0.03fF
C2751 _511_/a_93_21# _511_/a_346_47# 0.05fF
C2752 _529_/a_109_297# _531_/C 0.13fF
C2753 _548_/a_226_297# _530_/X 0.01fF
C2754 _561_/A _628_/Y 0.11fF
C2755 _567_/B _475_/A 0.02fF
C2756 _566_/A _386_/A 0.02fF
C2757 _626_/a_109_47# _626_/a_397_297# 0.05fF
C2758 _328_/A _314_/X 1.05fF
C2759 _567_/B _488_/X 0.41fF
C2760 _389_/a_27_47# VPWR 0.57fF
C2761 _603_/Y _604_/a_80_21# 0.30fF
C2762 _444_/A _442_/a_303_47# 0.06fF
C2763 _474_/A _472_/B 0.09fF
C2764 _569_/A _583_/X 0.01fF
C2765 _458_/X _460_/a_76_199# 0.07fF
C2766 B[7] _628_/Y 3.99fF
C2767 _343_/a_76_199# _343_/a_226_47# 0.49fF
C2768 _614_/a_226_47# _588_/A 0.14fF
C2769 _547_/a_222_93# _542_/D 0.00fF
C2770 _569_/Y _622_/C 0.03fF
C2771 _419_/a_76_199# VPWR 0.49fF
C2772 _428_/a_81_21# VPWR 0.44fF
C2773 _383_/X _442_/A 0.35fF
C2774 _554_/X _524_/a_78_199# 0.01fF
C2775 _521_/a_78_199# _483_/X 0.26fF
C2776 _583_/a_76_199# _583_/a_226_47# 0.49fF
C2777 _628_/a_300_47# _621_/X 0.32fF
C2778 _375_/a_544_297# VPWR 0.01fF
C2779 _420_/X _475_/A 0.19fF
C2780 _447_/a_68_297# _542_/A 0.01fF
C2781 _455_/X _485_/A 0.05fF
C2782 _406_/a_113_47# _433_/Y 0.05fF
C2783 VPWR _508_/a_323_297# 0.02fF
C2784 _495_/a_76_199# VPWR 0.71fF
C2785 VPWR _316_/a_558_47# 0.24fF
C2786 VPWR _363_/a_68_297# 0.34fF
C2787 _503_/a_664_47# _471_/A 0.20fF
C2788 _629_/B _432_/B 0.22fF
C2789 _513_/A _565_/a_80_21# 0.21fF
C2790 _555_/a_215_297# _555_/a_382_47# 0.03fF
C2791 _580_/A _578_/a_78_199# 0.06fF
C2792 _577_/a_226_47# _550_/X 0.01fF
C2793 _475_/a_68_297# _390_/B 0.08fF
C2794 _378_/a_62_47# _378_/a_381_47# 0.08fF
C2795 _561_/A _452_/X 0.75fF
C2796 _488_/a_76_199# _559_/a_77_199# 0.01fF
C2797 _365_/a_299_297# _371_/B 0.13fF
C2798 _585_/B _485_/D 0.26fF
C2799 _436_/A _331_/a_27_47# 0.38fF
C2800 _546_/a_226_47# _546_/X 0.05fF
C2801 _583_/X _627_/D 0.30fF
C2802 _516_/A _376_/X 0.01fF
C2803 _456_/a_76_199# _446_/X 0.01fF
C2804 _633_/Y _472_/Y 0.21fF
C2805 _580_/A _606_/A 0.18fF
C2806 _342_/X _328_/A 0.20fF
C2807 B[1] _380_/A 0.89fF
C2808 B[7] _452_/X 0.31fF
C2809 _475_/A _411_/A 0.48fF
C2810 _627_/D _622_/X 0.27fF
C2811 _398_/a_76_199# _398_/a_489_413# 0.12fF
C2812 _634_/Y _635_/a_27_413# 0.23fF
C2813 _365_/a_81_21# VPWR 0.42fF
C2814 _611_/X _442_/D 0.02fF
C2815 _619_/Y _607_/a_78_199# 0.01fF
C2816 _563_/a_27_297# VPWR 0.38fF
C2817 input7/a_27_47# _521_/a_215_47# 0.01fF
C2818 A[6] _521_/a_78_199# 0.01fF
C2819 _350_/X _397_/X 0.61fF
C2820 _338_/X _369_/a_226_47# 0.02fF
C2821 _352_/a_222_93# _352_/X 0.05fF
C2822 _352_/a_448_47# _328_/X 0.23fF
C2823 _411_/a_68_297# VPWR 0.27fF
C2824 _463_/a_76_199# _463_/a_226_47# 0.49fF
C2825 _585_/B _483_/X 0.84fF
C2826 _598_/a_68_297# _574_/X 0.00fF
C2827 B[1] _384_/a_226_47# 0.06fF
C2828 _539_/X _469_/X 0.10fF
C2829 _376_/a_68_297# _376_/a_150_297# 0.02fF
C2830 _454_/X _511_/a_250_297# 0.26fF
C2831 _357_/a_27_47# VPWR 0.34fF
C2832 _569_/A _589_/a_489_413# 0.09fF
C2833 _530_/X _547_/a_79_199# 0.17fF
C2834 A[3] _542_/A 0.36fF
C2835 _384_/X _396_/a_93_21# 0.01fF
C2836 _611_/X _588_/Y 1.44fF
C2837 _564_/a_219_297# _627_/a_27_297# 0.01fF
C2838 _613_/X _588_/A 0.77fF
C2839 _582_/a_27_47# _557_/Y 0.16fF
C2840 _517_/a_68_297# _517_/a_150_297# 0.02fF
C2841 input4/a_27_47# A[3] 0.41fF
C2842 _445_/A _519_/A 0.24fF
C2843 _491_/X _523_/X 0.24fF
C2844 _613_/a_77_199# _612_/Y 0.14fF
C2845 _331_/a_27_47# _350_/X 0.02fF
C2846 input3/a_62_47# A[2] 0.51fF
C2847 input3/a_664_47# input3/a_841_47# 0.29fF
C2848 _499_/a_81_21# _531_/A 0.25fF
C2849 _567_/Y _503_/A 0.15fF
C2850 _567_/B _511_/X 0.03fF
C2851 _468_/X VPWR 6.45fF
C2852 _454_/X _447_/B 0.03fF
C2853 _380_/A _383_/X 0.46fF
C2854 _635_/a_300_297# VPWR 0.55fF
C2855 _361_/X _363_/B 0.01fF
C2856 output31/a_27_47# _427_/Y 0.00fF
C2857 B[0] _503_/A 0.05fF
C2858 _542_/B _381_/B 0.21fF
C2859 _623_/a_489_413# _622_/X 0.14fF
C2860 _488_/a_489_413# _535_/Y 0.00fF
C2861 _386_/a_381_47# _386_/a_558_47# 0.32fF
C2862 _347_/A _313_/A 0.18fF
C2863 _567_/B _390_/B 0.03fF
C2864 _351_/A _371_/B 0.03fF
C2865 _590_/A _622_/a_29_53# 0.03fF
C2866 _420_/X _391_/a_150_297# 0.01fF
C2867 _516_/A M[9] 0.01fF
C2868 _585_/B A[6] 0.61fF
C2869 _410_/B _340_/A 0.20fF
C2870 M[7] _558_/a_77_199# 0.05fF
C2871 _567_/B _493_/X 0.29fF
C2872 _491_/a_76_199# _491_/a_226_297# 0.01fF
C2873 _491_/a_226_47# _491_/a_489_413# 0.02fF
C2874 _594_/a_27_297# _573_/Y 0.44fF
C2875 VPWR _628_/Y 3.82fF
C2876 _486_/a_68_297# _486_/X 0.27fF
C2877 _611_/a_109_47# _591_/A 0.05fF
C2878 _583_/X _579_/a_59_75# 0.06fF
C2879 _315_/a_161_47# _519_/C 0.02fF
C2880 _629_/X M[5] 0.14fF
C2881 _536_/Y _535_/Y 0.44fF
C2882 _530_/a_226_47# _531_/B 0.25fF
C2883 _417_/A _351_/X 0.08fF
C2884 _383_/X _384_/a_226_47# 0.53fF
C2885 _563_/B _485_/D 0.16fF
C2886 _563_/A _486_/A 0.39fF
C2887 _327_/a_215_47# _510_/A 0.16fF
C2888 _631_/Y VPWR 12.21fF
C2889 _429_/a_489_413# _398_/X 0.14fF
C2890 _412_/X _421_/a_226_47# 0.01fF
C2891 _614_/a_76_199# _611_/X 0.21fF
C2892 _360_/a_489_413# _359_/X 0.14fF
C2893 _533_/X _510_/A 0.01fF
C2894 _410_/a_27_47# _442_/B 0.01fF
C2895 _390_/B _468_/a_78_199# 0.17fF
C2896 _575_/a_78_199# _575_/a_292_297# 0.03fF
C2897 VPWR _621_/a_292_297# 0.01fF
C2898 _510_/a_68_297# _472_/Y 0.05fF
C2899 _597_/a_78_199# _597_/a_215_47# 0.26fF
C2900 _510_/A _473_/a_227_47# 0.02fF
C2901 _410_/a_27_47# _542_/B 0.46fF
C2902 _487_/X _469_/X 0.05fF
C2903 _569_/Y _587_/A 0.03fF
C2904 input12/a_558_47# _620_/X 0.01fF
C2905 _485_/A _547_/a_448_47# 0.07fF
C2906 _390_/D _563_/A 0.30fF
C2907 _336_/a_78_199# _314_/a_68_297# 0.00fF
C2908 _463_/a_76_199# _498_/A 0.01fF
C2909 _382_/X VPWR 1.77fF
C2910 _486_/a_68_297# _486_/a_150_297# 0.02fF
C2911 VPWR _397_/a_226_47# 0.16fF
C2912 _627_/C _586_/a_76_199# 0.14fF
C2913 _569_/Y _612_/A 0.26fF
C2914 _586_/S _433_/Y 0.12fF
C2915 _423_/X _631_/A 0.08fF
C2916 _627_/X _442_/D 0.76fF
C2917 _381_/C _484_/a_215_47# 0.12fF
C2918 _452_/X VPWR 2.17fF
C2919 _384_/X _397_/a_226_297# 0.05fF
C2920 _519_/a_111_297# _542_/A 0.01fF
C2921 _506_/A _480_/Y 0.99fF
C2922 _633_/Y _590_/B 0.03fF
C2923 _497_/B _463_/a_489_413# 0.01fF
C2924 _436_/A _384_/a_489_413# 0.02fF
C2925 _612_/Y _627_/A 0.08fF
C2926 _390_/B _411_/A 0.10fF
C2927 _390_/D _627_/A 0.10fF
C2928 _503_/a_381_47# VPWR 0.30fF
C2929 _626_/Y _525_/a_226_47# 0.10fF
C2930 _476_/a_250_297# _510_/A 0.00fF
C2931 _579_/a_59_75# _580_/a_68_297# 0.02fF
C2932 _506_/Y _533_/a_539_297# 0.02fF
C2933 _482_/a_68_297# _482_/X 0.27fF
C2934 A[6] _447_/X 0.13fF
C2935 VPWR _481_/a_27_47# 0.55fF
C2936 _569_/A _469_/A 0.36fF
C2937 _360_/a_76_199# _360_/X 0.22fF
C2938 _433_/Y _540_/X 0.04fF
C2939 _569_/Y _625_/Y 0.09fF
C2940 output24/a_27_47# VPWR 0.50fF
C2941 _505_/a_303_47# _482_/X 0.01fF
C2942 _544_/A _567_/Y 0.02fF
C2943 _390_/D _548_/X 0.47fF
C2944 _328_/B _420_/X 0.17fF
C2945 _506_/A _539_/A 0.02fF
C2946 VPWR _607_/a_215_47# 0.15fF
C2947 _544_/A B[0] 0.10fF
C2948 _417_/A _419_/X 1.00fF
C2949 _378_/a_841_47# _324_/a_664_47# 0.01fF
C2950 _533_/X _483_/X 0.27fF
C2951 _497_/A _527_/Y 0.20fF
C2952 _413_/X _417_/A 0.01fF
C2953 _327_/a_215_47# _631_/A 0.24fF
C2954 _529_/Y _531_/B 1.44fF
C2955 _455_/X _383_/X 0.07fF
C2956 _417_/D _512_/a_493_297# 0.02fF
C2957 _461_/a_215_47# _423_/X 0.10fF
C2958 _563_/B A[6] 0.66fF
C2959 _563_/D _381_/B 0.36fF
C2960 _570_/A _469_/X 0.12fF
C2961 _455_/X _356_/a_215_47# 0.11fF
C2962 B[1] _397_/a_76_199# 0.02fF
C2963 _542_/B _542_/A 0.88fF
C2964 _565_/a_80_21# _561_/A 0.00fF
C2965 _490_/a_78_199# VPWR 0.60fF
C2966 _486_/B _486_/X 0.01fF
C2967 _584_/A _530_/X 0.05fF
C2968 _457_/a_76_199# VPWR 0.49fF
C2969 _575_/a_215_47# _546_/X 0.11fF
C2970 _324_/a_664_47# _367_/C 0.12fF
C2971 _347_/A _512_/a_493_297# 0.08fF
C2972 _380_/a_27_47# _485_/A 0.13fF
C2973 _559_/X _575_/X 0.04fF
C2974 _606_/Y _607_/a_215_47# 0.11fF
C2975 _550_/X _521_/X 0.01fF
C2976 _335_/a_558_47# VPWR 0.23fF
C2977 _474_/A _446_/X 0.42fF
C2978 _355_/A VPWR 1.14fF
C2979 _626_/Y _591_/A 0.17fF
C2980 _513_/A _486_/B 0.07fF
C2981 _476_/X _633_/Y 0.51fF
C2982 _358_/a_27_47# _359_/B 0.20fF
C2983 input5/a_664_47# _431_/a_76_199# 0.00fF
C2984 _534_/a_80_21# _386_/A 0.27fF
C2985 B[6] _558_/X 0.10fF
C2986 _611_/a_27_297# _622_/C 0.11fF
C2987 _412_/X _419_/X 0.19fF
C2988 _451_/a_27_47# _563_/B 0.22fF
C2989 _567_/Y _566_/Y 0.62fF
C2990 _551_/a_76_199# _552_/a_489_413# 0.02fF
C2991 _551_/a_226_47# _552_/a_226_47# 0.00fF
C2992 _551_/a_489_413# _552_/a_76_199# 0.02fF
C2993 _362_/a_76_199# _351_/a_219_297# 0.01fF
C2994 _526_/a_76_199# VPWR 0.51fF
C2995 _332_/X _366_/a_489_413# 0.07fF
C2996 VPWR _624_/a_489_47# 0.03fF
C2997 _513_/a_27_47# _534_/a_209_297# 0.02fF
C2998 _603_/a_27_47# _554_/B 0.01fF
C2999 _603_/Y _555_/a_215_297# 0.16fF
C3000 _567_/Y _567_/a_109_297# 0.02fF
C3001 _328_/B _328_/X 0.01fF
C3002 _379_/a_292_297# VPWR 0.01fF
C3003 _360_/X _353_/X 0.03fF
C3004 _574_/X _616_/A 0.03fF
C3005 _561_/a_27_47# _454_/a_76_199# 0.01fF
C3006 _561_/A _447_/B 0.60fF
C3007 _575_/X _616_/B 0.21fF
C3008 _315_/a_161_47# _381_/C 0.56fF
C3009 _489_/a_226_297# _489_/a_76_199# 0.01fF
C3010 _625_/a_27_47# _606_/A 0.17fF
C3011 _322_/A _346_/A 0.14fF
C3012 _424_/X _390_/B 0.57fF
C3013 _382_/B _420_/a_222_93# 0.25fF
C3014 _591_/Y _599_/Y 1.07fF
C3015 _383_/X _397_/a_76_199# 0.01fF
C3016 _520_/a_226_47# VPWR 0.08fF
C3017 _518_/a_250_297# _381_/B 0.04fF
C3018 _510_/A _472_/a_109_297# 0.01fF
C3019 _380_/A _547_/X 0.03fF
C3020 _539_/A _515_/A 0.16fF
C3021 _516_/A _515_/A 0.39fF
C3022 _406_/A _458_/a_78_199# 0.12fF
C3023 _461_/X _462_/a_489_413# 0.16fF
C3024 _383_/X _452_/A 0.10fF
C3025 _503_/A _572_/A 0.63fF
C3026 _492_/X _504_/X 0.09fF
C3027 _574_/X _572_/A 0.02fF
C3028 B[7] _585_/a_109_297# 0.02fF
C3029 B[1] _335_/a_381_47# 0.14fF
C3030 _356_/a_215_47# _452_/A 0.03fF
C3031 _497_/A _531_/A 0.15fF
C3032 _386_/A _530_/X 0.10fF
C3033 input12/a_558_47# VPWR 0.22fF
C3034 _341_/a_27_47# _458_/X 0.07fF
C3035 _421_/a_226_47# _631_/B 0.07fF
C3036 _456_/X _457_/X 0.01fF
C3037 _615_/a_215_47# _573_/A 0.24fF
C3038 _330_/A _363_/B 0.03fF
C3039 _327_/a_78_199# _327_/a_292_297# 0.03fF
C3040 _587_/A _507_/Y 0.20fF
C3041 _541_/a_292_297# VPWR 0.02fF
C3042 _630_/a_226_47# _630_/X 0.05fF
C3043 _324_/a_62_47# _324_/a_558_47# 0.03fF
C3044 _543_/B _587_/A 0.11fF
C3045 _550_/X _550_/a_215_47# 0.01fF
C3046 _422_/a_489_413# _412_/X 0.07fF
C3047 _436_/A _503_/A 0.03fF
C3048 _549_/X _576_/X 0.15fF
C3049 _387_/a_292_297# _633_/Y 0.02fF
C3050 _432_/A _426_/A 0.08fF
C3051 _539_/A _535_/Y 0.10fF
C3052 _475_/X _475_/A 0.42fF
C3053 _487_/X _488_/a_226_47# 0.58fF
C3054 M[12] _442_/D 0.31fF
C3055 _546_/X _570_/A 0.18fF
C3056 _390_/B _426_/A 0.03fF
C3057 _478_/A _483_/a_250_297# 0.01fF
C3058 _504_/a_77_199# _468_/a_78_199# 0.01fF
C3059 _578_/a_78_199# _551_/X 0.27fF
C3060 _563_/A _563_/a_27_297# 0.34fF
C3061 _424_/a_226_47# _422_/X 0.22fF
C3062 _424_/a_489_413# _423_/X 0.14fF
C3063 _473_/a_77_199# _473_/a_539_297# 0.06fF
C3064 _563_/D _542_/A 0.03fF
C3065 _583_/X _448_/A 0.01fF
C3066 _534_/a_80_21# _386_/X 0.03fF
C3067 _504_/a_227_47# _510_/A 0.20fF
C3068 _362_/a_226_297# _351_/X 0.05fF
C3069 _554_/A _554_/B 1.23fF
C3070 _503_/A _542_/D 0.05fF
C3071 _313_/a_27_47# VPWR 0.54fF
C3072 _417_/A _338_/X 0.35fF
C3073 _608_/a_78_199# _609_/a_209_297# 0.02fF
C3074 _570_/a_150_297# _570_/A 0.01fF
C3075 _347_/A _408_/B 0.02fF
C3076 _363_/A _371_/A 0.03fF
C3077 _605_/a_209_297# _602_/Y 0.07fF
C3078 _543_/B _544_/a_558_47# 0.08fF
C3079 _408_/B _332_/X 0.20fF
C3080 _568_/a_539_297# _570_/B 0.08fF
C3081 _417_/D _488_/a_226_297# 0.02fF
C3082 _396_/a_346_47# _330_/A 0.05fF
C3083 _627_/C A[6] 0.27fF
C3084 _538_/Y _587_/A 0.15fF
C3085 _417_/D _472_/B 0.56fF
C3086 _609_/a_209_297# _542_/D 0.18fF
C3087 _442_/a_27_47# _316_/a_664_47# 0.01fF
C3088 _565_/a_80_21# VPWR 0.35fF
C3089 _500_/a_78_199# VPWR 0.78fF
C3090 _620_/a_226_297# _618_/A 0.02fF
C3091 _627_/A _357_/a_27_47# 0.09fF
C3092 _604_/a_80_21# _558_/a_77_199# 0.01fF
C3093 _628_/a_382_297# _628_/a_734_297# 0.02fF
C3094 _518_/X _381_/B 0.62fF
C3095 _530_/a_226_47# _530_/a_489_413# 0.02fF
C3096 _530_/a_76_199# _530_/a_226_297# 0.01fF
C3097 _442_/a_27_47# _443_/B 0.21fF
C3098 _375_/X M[2] 0.12fF
C3099 _543_/B _514_/a_68_297# 0.00fF
C3100 _542_/a_303_47# _542_/C 0.09fF
C3101 _476_/a_93_21# _390_/B 0.18fF
C3102 _631_/a_109_297# VPWR 0.01fF
C3103 _545_/Y VPWR 2.59fF
C3104 _437_/a_448_47# VPWR 0.04fF
C3105 _445_/A _337_/A 0.06fF
C3106 _546_/X _535_/A 0.08fF
C3107 _384_/X _363_/A 0.04fF
C3108 _563_/D _512_/a_292_297# 0.08fF
C3109 _544_/A _418_/a_68_297# 0.02fF
C3110 _626_/Y _520_/X 0.20fF
C3111 _464_/A _497_/A 0.26fF
C3112 _390_/D _333_/a_27_47# 0.50fF
C3113 _351_/X _374_/a_215_47# 0.11fF
C3114 _347_/A _445_/a_68_297# 0.20fF
C3115 _545_/Y _544_/a_664_47# 0.01fF
C3116 _581_/a_27_93# _581_/a_206_47# 0.02fF
C3117 _594_/X _593_/Y 0.42fF
C3118 _511_/a_250_297# VPWR 0.74fF
C3119 _488_/a_226_47# _570_/A 0.01fF
C3120 _468_/X _627_/A 0.01fF
C3121 _529_/Y _498_/A 0.24fF
C3122 _538_/A _469_/A 0.23fF
C3123 _503_/A _478_/A 0.27fF
C3124 _583_/X _601_/A 0.47fF
C3125 _359_/A _481_/A 0.49fF
C3126 _605_/a_80_21# _582_/a_27_47# 0.03fF
C3127 _630_/a_226_297# _432_/B 0.02fF
C3128 _326_/A VPWR 2.03fF
C3129 _585_/B _590_/B 0.16fF
C3130 _542_/A _489_/a_226_47# 0.00fF
C3131 B[1] _350_/a_27_297# 0.04fF
C3132 _419_/X _631_/B 2.67fF
C3133 _550_/X _580_/B 0.01fF
C3134 _583_/a_76_199# VPWR 0.50fF
C3135 _375_/X _332_/X 0.03fF
C3136 _417_/a_303_47# _519_/A 0.03fF
C3137 _337_/a_68_297# _338_/a_222_93# 0.00fF
C3138 A[4] VPWR 0.44fF
C3139 _473_/a_227_47# _472_/Y 0.05fF
C3140 VPWR _447_/B 2.65fF
C3141 _575_/X _530_/X 0.71fF
C3142 _475_/A _367_/a_27_297# 0.41fF
C3143 _419_/a_76_199# _419_/a_489_413# 0.12fF
C3144 _395_/a_68_297# _395_/a_150_297# 0.02fF
C3145 _587_/A _486_/X 0.32fF
C3146 _593_/A _591_/A 0.21fF
C3147 _455_/a_79_199# _419_/a_76_199# 0.00fF
C3148 _585_/a_109_297# VPWR 0.01fF
C3149 _619_/Y _606_/A 0.25fF
C3150 _595_/X _575_/a_78_199# 0.02fF
C3151 _456_/a_489_413# _456_/X 0.09fF
C3152 _540_/a_93_21# _469_/X 0.26fF
C3153 _493_/a_78_199# _457_/X 0.01fF
C3154 _532_/a_489_47# _527_/Y 0.16fF
C3155 _350_/C _481_/A 0.38fF
C3156 _627_/A _631_/Y 0.03fF
C3157 _613_/a_227_297# _627_/D 0.01fF
C3158 _542_/D _627_/a_205_297# 0.01fF
C3159 input10/a_27_47# _363_/A 0.14fF
C3160 _627_/X _627_/a_27_297# 0.20fF
C3161 _487_/a_215_47# _452_/X 0.10fF
C3162 _544_/A _542_/D 1.43fF
C3163 _633_/Y _350_/C 0.14fF
C3164 _633_/a_74_47# _367_/a_27_297# 0.00fF
C3165 _419_/X _411_/X 0.25fF
C3166 _634_/a_27_413# _337_/X 0.01fF
C3167 output19/a_27_47# _583_/X 0.40fF
C3168 VPWR _376_/a_68_297# 0.32fF
C3169 _561_/A _486_/B 0.01fF
C3170 _538_/A _559_/a_227_47# 0.14fF
C3171 _538_/Y _559_/a_323_297# 0.03fF
C3172 _316_/a_558_47# _316_/a_841_47# 0.07fF
C3173 _443_/B _316_/a_664_47# 0.01fF
C3174 _476_/a_93_21# _471_/A 0.01fF
C3175 _476_/a_256_47# _471_/Y 0.03fF
C3176 _506_/Y _585_/B 0.97fF
C3177 _495_/a_76_199# _495_/a_489_413# 0.12fF
C3178 _527_/B _527_/Y 1.04fF
C3179 _530_/a_489_413# _529_/Y 0.14fF
C3180 _520_/X _381_/B 0.43fF
C3181 _516_/A _382_/B 0.20fF
C3182 _475_/X _390_/B 1.34fF
C3183 _436_/A _391_/B 0.04fF
C3184 _566_/A _515_/A 0.03fF
C3185 _444_/Y _411_/A 0.08fF
C3186 _595_/a_77_199# _595_/a_539_297# 0.06fF
C3187 _622_/C _627_/B 0.13fF
C3188 _546_/a_76_199# _588_/A 0.01fF
C3189 _469_/A _488_/X 0.31fF
C3190 _386_/a_381_47# VPWR 0.30fF
C3191 _628_/a_382_297# B[7] 0.13fF
C3192 _362_/a_76_199# _351_/A 0.01fF
C3193 _481_/A _367_/C 0.04fF
C3194 _561_/A _418_/X 0.13fF
C3195 _408_/X _394_/a_558_47# 0.02fF
C3196 _491_/a_226_47# VPWR 0.12fF
C3197 _543_/Y _546_/a_489_413# 0.07fF
C3198 _445_/a_68_297# _445_/a_150_297# 0.02fF
C3199 _587_/A _454_/X 0.03fF
C3200 _566_/A _546_/a_76_199# 0.17fF
C3201 _515_/Y _546_/a_489_413# 0.02fF
C3202 _633_/Y _367_/C 0.20fF
C3203 _503_/a_381_47# _627_/A 0.79fF
C3204 _633_/a_265_297# VPWR 0.01fF
C3205 _382_/A _417_/A 0.41fF
C3206 _361_/a_226_47# _374_/X 0.02fF
C3207 A[3] _539_/A 0.98fF
C3208 _442_/A _481_/A 0.47fF
C3209 _386_/A _514_/B 0.68fF
C3210 _597_/a_292_297# VPWR 0.01fF
C3211 _351_/A _351_/a_219_297# 0.32fF
C3212 _493_/a_78_199# _459_/X 0.42fF
C3213 VPWR _486_/a_68_297# 0.34fF
C3214 _519_/A _484_/a_78_199# 0.39fF
C3215 _534_/a_80_21# _534_/a_209_47# 0.04fF
C3216 _448_/a_68_297# _448_/a_150_297# 0.02fF
C3217 _389_/a_27_47# _333_/a_27_47# 0.01fF
C3218 _471_/Y _478_/A 0.36fF
C3219 _556_/Y _582_/Y 0.00fF
C3220 _352_/X B[5] 0.03fF
C3221 B[7] _549_/a_226_297# 0.02fF
C3222 _569_/A _547_/X 0.02fF
C3223 _479_/B _482_/X 0.21fF
C3224 _360_/a_556_47# VPWR 0.00fF
C3225 VPWR _343_/X 0.43fF
C3226 _433_/Y _540_/a_346_47# 0.05fF
C3227 _313_/A _584_/A 0.35fF
C3228 _599_/A _597_/a_78_199# 0.00fF
C3229 _604_/X _558_/a_227_47# 0.01fF
C3230 _494_/a_489_413# VPWR 0.39fF
C3231 _618_/Y _620_/X 0.03fF
C3232 B[7] _622_/C 0.66fF
C3233 _455_/a_222_93# _455_/X 0.05fF
C3234 _485_/A _390_/B 1.03fF
C3235 _469_/a_381_47# _584_/A 0.10fF
C3236 B[1] _475_/A 0.20fF
C3237 _586_/a_76_199# _469_/X 0.01fF
C3238 _485_/a_109_47# _542_/D 0.02fF
C3239 _553_/a_292_297# _525_/X 0.04fF
C3240 _456_/X _504_/X 0.34fF
C3241 _386_/A _385_/a_381_47# 0.61fF
C3242 _491_/a_489_413# _490_/X 0.17fF
C3243 _553_/a_78_199# _524_/X 0.13fF
C3244 _563_/a_27_297# _563_/a_205_297# 0.01fF
C3245 _329_/a_76_199# _328_/X 0.22fF
C3246 _488_/X _489_/a_76_199# 0.14fF
C3247 _475_/X _471_/A 0.03fF
C3248 _561_/a_27_47# _627_/C 0.22fF
C3249 _495_/a_489_413# _468_/X 0.16fF
C3250 _495_/a_226_47# _494_/X 0.53fF
C3251 B[2] _485_/D 0.31fF
C3252 B[1] _633_/a_74_47# 0.23fF
C3253 _426_/A _371_/A 0.56fF
C3254 M[8] _558_/X 0.14fF
C3255 _412_/X _437_/a_222_93# 0.00fF
C3256 _595_/a_227_47# _570_/X 0.09fF
C3257 _412_/a_226_297# _408_/X 0.02fF
C3258 _467_/Y _467_/a_109_47# 0.47fF
C3259 _338_/X _631_/B 0.15fF
C3260 _547_/a_448_47# _547_/X 0.01fF
C3261 _457_/X _406_/Y 0.02fF
C3262 _633_/Y _610_/A 0.17fF
C3263 output31/a_27_47# _427_/A 0.01fF
C3264 _458_/X VPWR 2.29fF
C3265 _408_/B _336_/a_78_199# 0.36fF
C3266 _557_/A B[6] 0.05fF
C3267 _476_/a_93_21# _504_/a_77_199# 0.08fF
C3268 _349_/a_493_297# _419_/X 0.02fF
C3269 _472_/a_109_297# _472_/Y 0.02fF
C3270 _573_/A _572_/A 0.47fF
C3271 _335_/a_841_47# _632_/a_215_47# 0.02fF
C3272 VPWR _522_/X 0.70fF
C3273 _568_/a_227_47# _469_/X 0.10fF
C3274 _431_/a_76_199# _431_/a_489_413# 0.12fF
C3275 _327_/a_78_199# VPWR 0.06fF
C3276 _461_/a_78_199# _461_/X 0.21fF
C3277 _416_/a_78_199# _448_/B 0.01fF
C3278 _469_/A _511_/X 0.01fF
C3279 _520_/X _542_/A 0.23fF
C3280 _578_/a_215_47# VPWR 0.05fF
C3281 _500_/a_78_199# _531_/C 0.21fF
C3282 _590_/A _593_/A 0.15fF
C3283 _380_/A _481_/A 1.81fF
C3284 _570_/B _503_/A 0.50fF
C3285 _473_/a_227_297# VPWR 0.01fF
C3286 _626_/Y _574_/X 0.20fF
C3287 _520_/X input4/a_27_47# 0.07fF
C3288 _383_/X _475_/A 0.51fF
C3289 _542_/B _480_/Y 0.12fF
C3290 _380_/A _633_/Y 0.03fF
C3291 _517_/a_68_297# _584_/A 0.30fF
C3292 _417_/A _631_/A 0.59fF
C3293 _448_/B M[9] 0.22fF
C3294 _417_/D _517_/X 0.36fF
C3295 _329_/a_76_199# _329_/X 0.24fF
C3296 _360_/X _361_/X 0.84fF
C3297 VPWR _624_/X 1.70fF
C3298 VPWR _486_/B 1.18fF
C3299 _455_/a_222_93# _452_/A 0.13fF
C3300 _337_/B _332_/X 0.12fF
C3301 _411_/B _437_/a_79_199# 0.22fF
C3302 _533_/X _506_/Y 0.01fF
C3303 _628_/a_382_297# VPWR 0.39fF
C3304 VPWR output18/a_27_47# 0.63fF
C3305 _441_/a_78_199# _346_/A 0.15fF
C3306 _347_/A _517_/X 0.10fF
C3307 _523_/X _631_/Y 0.39fF
C3308 _603_/Y _631_/Y 0.04fF
C3309 _439_/X _468_/a_292_297# 0.08fF
C3310 _581_/a_27_93# VPWR 0.31fF
C3311 _510_/A _469_/X 0.24fF
C3312 _459_/X _406_/Y 0.02fF
C3313 _527_/A _557_/Y 0.00fF
C3314 _630_/X _397_/X 0.34fF
C3315 _520_/a_76_199# _547_/X 0.00fF
C3316 _519_/X _547_/a_222_93# 0.36fF
C3317 _370_/A _635_/a_300_297# 0.12fF
C3318 _530_/X M[9] 0.04fF
C3319 _628_/a_28_47# _623_/X 0.31fF
C3320 _599_/A _601_/A 0.09fF
C3321 _461_/a_78_199# _407_/a_27_47# 0.04fF
C3322 _418_/X VPWR 1.41fF
C3323 _586_/S _564_/A 0.52fF
C3324 _342_/X _343_/X 1.78fF
C3325 _445_/A VPWR 2.89fF
C3326 _468_/a_215_47# _437_/X 0.11fF
C3327 _589_/a_76_199# _589_/a_226_47# 0.49fF
C3328 _626_/Y _427_/A 0.03fF
C3329 _579_/X _554_/B 0.01fF
C3330 _375_/X _336_/a_78_199# 0.13fF
C3331 _406_/Y _503_/A 0.02fF
C3332 _635_/Y VPWR 0.43fF
C3333 _542_/B _539_/A 0.03fF
C3334 _567_/Y _539_/X 0.01fF
C3335 _467_/Y _527_/A 0.36fF
C3336 _516_/A _542_/B 0.03fF
C3337 _587_/A _537_/a_77_199# 0.24fF
C3338 _395_/a_68_297# VPWR 0.30fF
C3339 _453_/a_346_47# _542_/D 0.06fF
C3340 _559_/X _535_/Y 0.01fF
C3341 _571_/a_93_21# _571_/a_250_297# 0.50fF
C3342 _433_/Y _507_/Y 0.03fF
C3343 _588_/A A[3] 0.07fF
C3344 B[0] _539_/X 0.11fF
C3345 _485_/D _469_/X 0.03fF
C3346 input3/a_381_47# _485_/D 0.12fF
C3347 _626_/Y _549_/a_76_199# 0.08fF
C3348 _427_/A _467_/a_109_47# 0.02fF
C3349 VPWR _350_/B 2.32fF
C3350 _466_/X _467_/a_397_297# 0.13fF
C3351 _475_/X _504_/a_77_199# 0.39fF
C3352 VPWR _622_/C 6.65fF
C3353 _566_/A A[3] 0.03fF
C3354 _612_/A _620_/X 0.04fF
C3355 _542_/B _478_/a_303_47# 0.03fF
C3356 _563_/D _340_/a_27_47# 0.32fF
C3357 _560_/a_27_47# _563_/B 0.45fF
C3358 _469_/A _595_/a_77_199# 0.08fF
C3359 _567_/B _390_/D 0.08fF
C3360 _629_/A _630_/a_226_47# 0.06fF
C3361 _625_/Y _627_/B 0.04fF
C3362 B[1] _390_/B 0.05fF
C3363 _448_/a_68_297# VPWR 0.32fF
C3364 _503_/A _381_/B 0.05fF
C3365 _627_/C _590_/B 0.48fF
C3366 _476_/X _476_/a_250_297# 0.03fF
C3367 _618_/Y VPWR 1.78fF
C3368 _474_/Y _478_/A 0.04fF
C3369 _519_/X _518_/X 1.27fF
C3370 B[7] _612_/A 0.11fF
C3371 _487_/X _479_/B 0.06fF
C3372 _469_/X _483_/X 0.05fF
C3373 _627_/A _545_/Y 0.32fF
C3374 _397_/X _363_/B 0.03fF
C3375 _625_/Y _620_/X 0.28fF
C3376 _611_/a_109_47# _591_/Y 0.02fF
C3377 _359_/X _359_/A 0.82fF
C3378 _538_/Y _433_/Y 0.70fF
C3379 _424_/a_226_47# _406_/Y 0.00fF
C3380 _378_/A _519_/A 0.28fF
C3381 _459_/a_489_413# _457_/X 0.07fF
C3382 _563_/A _326_/A 0.74fF
C3383 B[2] _598_/B 0.03fF
C3384 _506_/Y _509_/Y 0.23fF
C3385 _606_/Y _618_/Y 0.33fF
C3386 _619_/a_27_47# _619_/Y 0.11fF
C3387 _455_/X _481_/A 0.07fF
C3388 _350_/X B[5] 0.27fF
C3389 _440_/a_556_47# _458_/X 0.02fF
C3390 _417_/D _442_/D 0.05fF
C3391 _424_/X _406_/B 0.01fF
C3392 _611_/a_109_297# _590_/B 0.00fF
C3393 _410_/C _472_/B 0.28fF
C3394 _589_/a_226_47# _612_/A 0.31fF
C3395 _433_/a_397_297# _433_/Y 0.20fF
C3396 _498_/Y _498_/A 0.34fF
C3397 _455_/X _633_/Y 0.11fF
C3398 _625_/Y B[7] 0.35fF
C3399 _429_/a_76_199# _371_/B 0.18fF
C3400 _543_/B _542_/a_27_47# 0.34fF
C3401 _604_/a_80_21# _604_/a_303_47# 0.04fF
C3402 A[6] _484_/a_215_47# 0.08fF
C3403 _444_/A _478_/A 0.24fF
C3404 _410_/C _445_/a_68_297# 0.16fF
C3405 _469_/a_62_47# _503_/A 0.07fF
C3406 _487_/X B[0] 0.50fF
C3407 _417_/D _417_/a_27_47# 0.23fF
C3408 _504_/a_77_199# _504_/a_539_297# 0.06fF
C3409 _582_/a_27_47# _556_/A 0.17fF
C3410 _390_/B _383_/X 0.57fF
C3411 _538_/Y _540_/X 1.19fF
C3412 _526_/a_76_199# _523_/X 0.01fF
C3413 _589_/a_76_199# VPWR 0.26fF
C3414 _603_/Y _526_/a_76_199# 0.13fF
C3415 _369_/a_489_413# B[5] 0.11fF
C3416 _376_/X _383_/a_226_47# 0.47fF
C3417 A[6] _469_/X 0.05fF
C3418 _534_/a_80_21# _515_/A 0.14fF
C3419 _594_/X _595_/X 2.86fF
C3420 _431_/X _466_/X 0.01fF
C3421 _626_/Y _504_/X 0.03fF
C3422 _585_/B _442_/A 0.41fF
C3423 _396_/X _397_/a_76_199# 0.24fF
C3424 _623_/X _589_/a_489_413# 0.11fF
C3425 _625_/Y _589_/a_226_47# 0.36fF
C3426 _328_/A _420_/X 0.13fF
C3427 _570_/B _566_/Y 0.34fF
C3428 _458_/a_78_199# _421_/X 0.29fF
C3429 _455_/X _490_/a_215_47# 0.14fF
C3430 _516_/A _563_/D 0.39fF
C3431 _504_/a_323_297# _587_/A 0.04fF
C3432 _436_/A _412_/a_226_297# 0.01fF
C3433 _563_/D _539_/A 0.30fF
C3434 _433_/Y _486_/X 0.07fF
C3435 _485_/D _546_/X 0.54fF
C3436 _408_/B _584_/A 1.32fF
C3437 _596_/a_76_199# _595_/X 0.21fF
C3438 _596_/a_226_47# _594_/X 0.22fF
C3439 _453_/X _519_/C 0.30fF
C3440 _437_/a_222_93# _411_/X 0.12fF
C3441 _573_/Y _574_/a_299_297# 0.05fF
C3442 VPWR _370_/B 0.84fF
C3443 _520_/X _523_/a_226_47# 0.01fF
C3444 _510_/A _411_/X 0.09fF
C3445 _542_/C _479_/B 0.66fF
C3446 _475_/A _438_/a_150_297# 0.01fF
C3447 _519_/X _520_/X 0.01fF
C3448 _544_/A _381_/B 0.35fF
C3449 VPWR _604_/a_209_297# 0.45fF
C3450 _425_/a_76_199# _425_/a_226_47# 0.49fF
C3451 _407_/Y _390_/B 0.25fF
C3452 _596_/a_76_199# _596_/a_226_47# 0.49fF
C3453 _504_/a_227_297# VPWR 0.01fF
C3454 _438_/X _468_/a_493_297# 0.12fF
C3455 _441_/a_215_47# VPWR 0.05fF
C3456 _516_/A _477_/a_292_297# 0.01fF
C3457 _503_/A _542_/A 0.05fF
C3458 _587_/A _439_/a_226_297# 0.02fF
C3459 _562_/a_215_47# _584_/A 0.16fF
C3460 _487_/a_78_199# _447_/X 0.33fF
C3461 _445_/X _445_/a_68_297# 0.27fF
C3462 _567_/Y _570_/A 0.68fF
C3463 _385_/a_62_47# _391_/B 0.12fF
C3464 _350_/C _409_/a_292_297# 0.07fF
C3465 B[1] _384_/a_226_297# 0.02fF
C3466 _503_/a_381_47# _503_/a_664_47# 0.09fF
C3467 _371_/B _373_/Y 0.01fF
C3468 _452_/A _481_/A 0.51fF
C3469 _338_/a_448_47# _338_/X 0.01fF
C3470 _328_/B _383_/X 0.29fF
C3471 _540_/X _486_/X 0.27fF
C3472 _508_/a_539_297# _507_/Y 0.02fF
C3473 _613_/X _613_/a_227_47# 0.04fF
C3474 _447_/X _367_/C 0.03fF
C3475 _536_/Y _520_/X 0.04fF
C3476 _534_/a_303_47# _381_/B 0.01fF
C3477 B[0] _570_/A 0.32fF
C3478 _530_/X _515_/A 0.52fF
C3479 _454_/X _433_/Y 0.03fF
C3480 _560_/a_27_47# _627_/C 0.07fF
C3481 _563_/a_27_297# _541_/a_215_47# 0.06fF
C3482 _566_/A _542_/B 0.07fF
C3483 _516_/a_27_47# _481_/a_27_47# 0.00fF
C3484 output25/a_27_47# _343_/X 0.01fF
C3485 _611_/a_27_297# _610_/Y 0.13fF
C3486 _591_/Y _626_/Y 0.03fF
C3487 _585_/B _610_/A 0.44fF
C3488 _440_/a_76_199# _478_/A 0.08fF
C3489 _631_/B _631_/A 1.22fF
C3490 _328_/A _328_/X 0.68fF
C3491 _587_/A VPWR 6.57fF
C3492 _425_/a_76_199# VPWR 0.57fF
C3493 _336_/a_78_199# _337_/B 0.21fF
C3494 VPWR _439_/a_489_413# 0.43fF
C3495 _371_/B VPWR 9.49fF
C3496 _542_/C B[0] 0.05fF
C3497 _360_/X _330_/A 0.12fF
C3498 _612_/A VPWR 3.68fF
C3499 _626_/Y _587_/a_27_47# 0.11fF
C3500 _453_/a_93_21# _453_/a_256_47# 0.03fF
C3501 _420_/a_222_93# _420_/a_448_47# 0.03fF
C3502 _326_/a_27_47# VPWR 0.53fF
C3503 _363_/A _363_/a_68_297# 0.34fF
C3504 _575_/X _575_/a_78_199# 0.21fF
C3505 _607_/X _607_/a_78_199# 0.21fF
C3506 _566_/Y _381_/B 0.71fF
C3507 _530_/X _535_/Y 0.10fF
C3508 _455_/X _413_/a_68_297# 0.20fF
C3509 _563_/B _367_/C 0.19fF
C3510 _605_/a_209_297# _557_/A 0.09fF
C3511 _348_/a_27_47# _475_/A 0.29fF
C3512 _518_/a_93_21# _517_/X 0.49fF
C3513 _447_/a_150_297# _542_/D 0.01fF
C3514 VPWR _361_/a_489_413# 0.39fF
C3515 _513_/A _542_/a_27_47# 0.01fF
C3516 _410_/a_27_47# _446_/a_93_21# 0.00fF
C3517 _544_/a_558_47# VPWR 0.22fF
C3518 _586_/S _451_/A 0.57fF
C3519 _625_/Y VPWR 2.99fF
C3520 _489_/a_226_47# _489_/X 0.05fF
C3521 _313_/A _395_/X 0.00fF
C3522 _493_/X _502_/a_78_199# 0.13fF
C3523 _519_/C _542_/D 0.40fF
C3524 _524_/a_78_199# _476_/X 0.31fF
C3525 _633_/Y _627_/D 0.12fF
C3526 _383_/X _384_/a_226_297# 0.01fF
C3527 _365_/a_81_21# _363_/A 0.17fF
C3528 _544_/a_381_47# _544_/a_841_47# 0.03fF
C3529 _544_/a_558_47# _544_/a_664_47# 0.60fF
C3530 _488_/a_76_199# _488_/X 0.22fF
C3531 _601_/Y VPWR 2.75fF
C3532 _382_/A _382_/a_68_297# 0.31fF
C3533 _327_/a_215_47# _367_/C 0.03fF
C3534 VPWR _514_/a_68_297# 0.41fF
C3535 _359_/X _380_/A 0.01fF
C3536 _503_/a_381_47# _475_/a_68_297# 0.02fF
C3537 _335_/a_381_47# _633_/Y 0.08fF
C3538 _342_/X _370_/B 0.03fF
C3539 _431_/a_226_47# _431_/X 0.05fF
C3540 _478_/A _430_/X 0.59fF
C3541 _613_/a_77_199# _622_/C 0.01fF
C3542 _487_/X _453_/X 0.01fF
C3543 _563_/A _486_/B 0.43fF
C3544 output19/a_27_47# output23/a_27_47# 0.01fF
C3545 _585_/B _508_/a_227_297# 0.03fF
C3546 _355_/A _478_/a_27_47# 0.05fF
C3547 _567_/B _468_/X 0.65fF
C3548 output31/a_27_47# _465_/a_27_297# 0.01fF
C3549 _490_/X VPWR 1.59fF
C3550 _577_/a_76_199# _577_/a_226_47# 0.49fF
C3551 _601_/Y _606_/Y 1.46fF
C3552 _351_/X _352_/X 0.17fF
C3553 _563_/D _340_/A 4.62fF
C3554 _496_/a_493_297# VPWR 0.01fF
C3555 _544_/A _542_/A 0.90fF
C3556 _554_/X _582_/a_27_47# 0.03fF
C3557 _561_/A _484_/a_78_199# 0.43fF
C3558 _514_/a_68_297# _514_/a_150_297# 0.02fF
C3559 _472_/Y _469_/X 0.04fF
C3560 _549_/X _551_/a_556_47# 0.02fF
C3561 _457_/a_76_199# _457_/a_489_413# 0.12fF
C3562 _404_/a_664_47# _503_/A 0.05fF
C3563 VPWR _559_/a_323_297# 0.01fF
C3564 _548_/a_76_199# _485_/D 0.07fF
C3565 _516_/A _518_/X 0.64fF
C3566 _408_/X _419_/X 0.62fF
C3567 _480_/A _479_/a_68_297# 0.27fF
C3568 _610_/A _616_/Y 0.44fF
C3569 _381_/C _453_/X 0.01fF
C3570 _375_/a_222_93# _359_/X 0.21fF
C3571 _378_/A _454_/X 0.03fF
C3572 _445_/A _563_/A 0.22fF
C3573 _411_/a_68_297# _411_/A 0.33fF
C3574 _335_/a_558_47# _335_/a_841_47# 0.07fF
C3575 _380_/A _334_/a_197_47# 0.03fF
C3576 _498_/A _466_/X 0.01fF
C3577 _439_/X _468_/a_215_47# 0.05fF
C3578 _440_/X _436_/X 0.03fF
C3579 _468_/X _468_/a_78_199# 0.21fF
C3580 _342_/X _371_/B 0.01fF
C3581 _329_/a_226_47# VPWR 0.07fF
C3582 _567_/B _631_/Y 0.03fF
C3583 _411_/B _446_/a_93_21# 0.04fF
C3584 _563_/A _350_/B 0.26fF
C3585 _386_/X _408_/B 0.01fF
C3586 _525_/a_76_199# _492_/a_76_199# 0.06fF
C3587 _469_/A _571_/a_584_47# 0.03fF
C3588 _482_/a_68_297# A[6] 0.15fF
C3589 _479_/a_68_297# _481_/A 0.10fF
C3590 A[1] _390_/B 0.04fF
C3591 _583_/X _612_/Y 0.03fF
C3592 _433_/Y _627_/B 2.54fF
C3593 _380_/A _563_/B 0.07fF
C3594 _382_/B _448_/B 0.26fF
C3595 _349_/a_292_297# _475_/A 0.08fF
C3596 _370_/a_68_297# output26/a_27_47# 0.01fF
C3597 _583_/X _390_/D 0.09fF
C3598 _526_/a_76_199# _526_/a_489_413# 0.12fF
C3599 _479_/A _518_/a_250_297# 0.02fF
C3600 _454_/X _316_/a_664_47# 0.12fF
C3601 _420_/X _631_/Y 0.03fF
C3602 _612_/Y _622_/X 0.01fF
C3603 _627_/A _622_/C 0.35fF
C3604 _586_/S _627_/B 1.45fF
C3605 _627_/A _595_/a_227_297# 0.03fF
C3606 _537_/a_77_199# _433_/Y 0.17fF
C3607 VPWR _466_/a_78_199# 0.60fF
C3608 input11/a_27_47# VPWR 0.51fF
C3609 _360_/X _442_/B 0.07fF
C3610 VPWR _361_/a_76_199# 0.46fF
C3611 _570_/X _469_/X 0.47fF
C3612 _569_/A _543_/Y 0.29fF
C3613 _361_/a_226_297# _361_/a_76_199# 0.01fF
C3614 _487_/X _542_/D 0.08fF
C3615 _404_/a_62_47# _622_/C 0.01fF
C3616 _390_/D _537_/a_227_297# 0.03fF
C3617 _471_/A _470_/a_209_297# 0.04fF
C3618 _387_/a_215_47# VPWR 0.05fF
C3619 _432_/A _629_/X 0.14fF
C3620 _585_/B _509_/A 0.03fF
C3621 _506_/Y _533_/a_77_199# 0.18fF
C3622 _356_/a_292_297# VPWR 0.01fF
C3623 input10/a_27_47# B[1] 0.41fF
C3624 _586_/a_505_21# _588_/A 0.01fF
C3625 _329_/a_226_47# _314_/X 0.31fF
C3626 _488_/a_489_413# _503_/A 0.01fF
C3627 _382_/X _420_/X 0.00fF
C3628 _514_/B _515_/A 0.01fF
C3629 _384_/X _383_/X 0.61fF
C3630 _631_/Y _411_/A 0.03fF
C3631 A[3] _530_/X 0.03fF
C3632 _515_/Y _518_/a_346_47# 0.02fF
C3633 _455_/X _359_/X 0.54fF
C3634 VPWR _399_/a_493_297# 0.01fF
C3635 _393_/A VPWR 2.56fF
C3636 _564_/a_219_297# _564_/a_27_53# 0.22fF
C3637 _516_/A _520_/X 0.40fF
C3638 _510_/X _533_/a_539_297# 0.02fF
C3639 _520_/X _539_/A 0.88fF
C3640 _375_/X _386_/X 0.02fF
C3641 _591_/Y _593_/A 1.53fF
C3642 B[7] _433_/Y 0.49fF
C3643 _381_/C _542_/D 2.48fF
C3644 _588_/a_109_297# _588_/Y 0.03fF
C3645 _428_/a_81_21# _426_/A 0.26fF
C3646 _588_/A _591_/A 0.47fF
C3647 _586_/S B[7] 0.04fF
C3648 _439_/X _504_/a_227_47# 0.01fF
C3649 _368_/B _634_/a_27_413# 0.03fF
C3650 _329_/a_226_47# _329_/a_489_413# 0.02fF
C3651 _329_/a_76_199# _329_/a_226_297# 0.01fF
C3652 _571_/a_256_47# _381_/B 0.01fF
C3653 B[0] _540_/a_93_21# 0.09fF
C3654 _436_/A _384_/a_76_199# 0.02fF
C3655 _584_/A _517_/X 0.06fF
C3656 _444_/A _410_/a_27_47# 0.16fF
C3657 _599_/Y _624_/a_585_369# 0.03fF
C3658 _529_/a_27_47# VPWR 0.03fF
C3659 _449_/A _453_/a_250_297# 0.05fF
C3660 _353_/X _375_/X 0.64fF
C3661 _627_/X _623_/a_76_199# 0.01fF
C3662 B[7] _540_/X 0.21fF
C3663 _370_/A _343_/X 0.45fF
C3664 _608_/X _610_/A 0.00fF
C3665 VPWR _484_/a_78_199# 0.58fF
C3666 _410_/B _472_/B 0.03fF
C3667 _340_/A _518_/X 0.40fF
C3668 _610_/Y _620_/X 0.10fF
C3669 _557_/A _531_/a_193_297# 0.14fF
C3670 _523_/X _522_/X 0.01fF
C3671 _573_/A _593_/A 0.67fF
C3672 _569_/A _585_/B 0.30fF
C3673 _442_/D _410_/C 1.37fF
C3674 _550_/X _552_/a_76_199# 0.01fF
C3675 _400_/a_80_21# VPWR 0.36fF
C3676 _551_/X _552_/a_226_47# 0.51fF
C3677 _533_/X _552_/a_489_413# 0.14fF
C3678 _417_/a_27_47# _311_/a_27_47# 0.01fF
C3679 _386_/a_62_47# _480_/A 0.00fF
C3680 _542_/C _542_/D 0.41fF
C3681 _626_/a_109_47# _624_/a_206_369# 0.04fF
C3682 _627_/C _610_/A 0.51fF
C3683 _419_/a_489_413# _418_/X 0.14fF
C3684 _385_/a_381_47# _385_/a_664_47# 0.09fF
C3685 input12/a_558_47# input12/a_841_47# 0.07fF
C3686 VPWR _555_/a_298_297# 0.42fF
C3687 _568_/a_77_199# _568_/a_539_297# 0.06fF
C3688 _455_/a_79_199# _418_/X 0.21fF
C3689 _561_/A _324_/a_381_47# 0.01fF
C3690 _528_/a_81_21# _527_/Y 0.33fF
C3691 _432_/A _432_/B 1.04fF
C3692 _537_/a_77_199# _537_/a_539_297# 0.06fF
C3693 _623_/X _613_/a_227_297# 0.01fF
C3694 _625_/Y _613_/a_77_199# 0.11fF
C3695 _570_/X _546_/X 0.34fF
C3696 _390_/D _485_/A 0.63fF
C3697 B[7] _610_/Y 0.35fF
C3698 _534_/a_80_21# _542_/B 0.11fF
C3699 _539_/a_68_297# _585_/B 0.06fF
C3700 _397_/X _398_/a_76_199# 0.25fF
C3701 _544_/A _519_/X 0.22fF
C3702 _516_/A _322_/A 0.46fF
C3703 _506_/Y _469_/X 0.03fF
C3704 M[8] _531_/A 0.77fF
C3705 _466_/a_78_199# _466_/a_292_297# 0.03fF
C3706 _475_/A _481_/A 0.47fF
C3707 _338_/X _344_/a_78_199# 0.13fF
C3708 _504_/a_227_297# _627_/A 0.01fF
C3709 _480_/Y _483_/a_250_297# 0.01fF
C3710 _380_/A _627_/C 0.06fF
C3711 _633_/Y _475_/A 5.42fF
C3712 _412_/a_76_199# _412_/a_489_413# 0.12fF
C3713 _378_/A _561_/A 3.24fF
C3714 _633_/Y _488_/X 0.52fF
C3715 _367_/a_109_297# _367_/C 0.04fF
C3716 _386_/A _517_/X 0.02fF
C3717 _408_/B _395_/X 0.31fF
C3718 _436_/A _419_/X 3.72fF
C3719 _611_/a_109_297# _610_/A 0.01fF
C3720 _544_/A _536_/Y 0.00fF
C3721 _563_/D _409_/a_215_47# 0.01fF
C3722 output25/a_27_47# _371_/B 0.10fF
C3723 _444_/A _411_/B 0.15fF
C3724 _455_/X _533_/X 0.29fF
C3725 _386_/X _458_/a_215_47# 0.13fF
C3726 _437_/X _631_/B 0.05fF
C3727 _373_/Y _433_/Y 0.01fF
C3728 _476_/X _469_/X 0.02fF
C3729 _356_/a_78_199# _356_/a_215_47# 0.26fF
C3730 _478_/A _508_/a_77_199# 0.09fF
C3731 _587_/A _627_/A 1.42fF
C3732 _633_/a_74_47# _633_/Y 0.32fF
C3733 _487_/a_493_297# VPWR 0.01fF
C3734 _533_/X _509_/A 0.04fF
C3735 _540_/a_346_47# _486_/X 0.02fF
C3736 _542_/C _478_/A 0.21fF
C3737 _419_/X _542_/D 1.86fF
C3738 _587_/A _438_/a_68_297# 0.00fF
C3739 _427_/Y _465_/X 0.01fF
C3740 _413_/X _542_/D 0.03fF
C3741 _381_/a_109_47# _381_/B 0.06fF
C3742 _485_/A _328_/A 0.03fF
C3743 _584_/A _442_/D 0.11fF
C3744 _520_/X _340_/A 0.03fF
C3745 VPWR _433_/Y 7.78fF
C3746 _542_/B _530_/X 0.05fF
C3747 _586_/S VPWR 4.52fF
C3748 _623_/X M[6] 0.07fF
C3749 _596_/a_76_199# _575_/X 0.01fF
C3750 _437_/X _411_/X 0.00fF
C3751 _510_/a_68_297# _510_/X 0.27fF
C3752 _568_/a_227_47# _567_/Y 0.05fF
C3753 _563_/B _452_/A 0.16fF
C3754 _390_/D _469_/A 0.05fF
C3755 _522_/a_76_199# _522_/a_226_47# 0.49fF
C3756 _571_/a_346_47# _469_/X 0.02fF
C3757 _355_/a_161_47# _355_/A 0.58fF
C3758 _625_/Y _627_/A 0.35fF
C3759 _362_/a_226_47# _371_/B 0.02fF
C3760 _417_/A _317_/a_27_47# 0.46fF
C3761 _635_/Y _370_/A 0.66fF
C3762 _590_/A _588_/A 0.24fF
C3763 _443_/B _446_/a_584_47# 0.03fF
C3764 M[8] _464_/A 0.17fF
C3765 _543_/B _565_/a_209_297# 0.03fF
C3766 _419_/X _350_/X 0.06fF
C3767 _628_/a_28_47# _628_/Y 0.27fF
C3768 _466_/a_215_47# _428_/X 0.24fF
C3769 _543_/A _545_/Y 0.03fF
C3770 VPWR _540_/X 5.21fF
C3771 _338_/a_79_199# _337_/A 0.39fF
C3772 _406_/B _405_/a_109_297# 0.02fF
C3773 _417_/a_27_47# _417_/a_109_47# 0.03fF
C3774 _362_/a_76_199# VPWR 0.48fF
C3775 _569_/A _572_/B 0.09fF
C3776 _573_/Y _547_/X 0.25fF
C3777 _492_/a_76_199# _492_/a_226_47# 0.49fF
C3778 _600_/a_114_47# _601_/A 0.01fF
C3779 _519_/A _376_/a_150_297# 0.02fF
C3780 _463_/a_489_413# _462_/X 0.21fF
C3781 _463_/a_226_297# _406_/Y 0.01fF
C3782 _444_/Y _470_/a_209_297# 0.09fF
C3783 _313_/A _391_/A 0.16fF
C3784 _565_/a_80_21# _565_/a_209_47# 0.04fF
C3785 _412_/X _406_/A 0.08fF
C3786 _351_/a_219_297# VPWR 0.24fF
C3787 _629_/X _371_/A 0.03fF
C3788 _386_/X _517_/X 0.41fF
C3789 input5/a_558_47# input5/a_664_47# 0.60fF
C3790 input5/a_381_47# input5/a_841_47# 0.03fF
C3791 _627_/D _616_/Y 0.02fF
C3792 _327_/a_215_47# _336_/a_215_47# 0.01fF
C3793 _577_/a_226_47# _576_/X 0.51fF
C3794 _577_/a_489_413# _559_/X 0.07fF
C3795 _503_/A _539_/A 1.72fF
C3796 _442_/a_27_47# VPWR 0.76fF
C3797 _616_/B _591_/A 0.14fF
C3798 _513_/A _520_/a_489_413# 0.09fF
C3799 _455_/X _509_/Y 0.16fF
C3800 _542_/a_27_47# VPWR 0.72fF
C3801 M[1] output24/a_27_47# 0.45fF
C3802 _633_/Y _511_/X 0.03fF
C3803 _513_/A _519_/A 0.13fF
C3804 _437_/a_222_93# _408_/X 0.03fF
C3805 _610_/Y VPWR 1.48fF
C3806 _512_/a_215_47# _514_/A 0.01fF
C3807 _406_/B _407_/Y 0.28fF
C3808 output27/a_27_47# _371_/A 0.00fF
C3809 _469_/a_381_47# _469_/a_664_47# 0.09fF
C3810 _574_/X _598_/A 0.11fF
C3811 _628_/Y _622_/X 0.26fF
C3812 VPWR _324_/a_381_47# 0.30fF
C3813 _509_/Y _509_/A 1.40fF
C3814 _322_/A _340_/A 0.44fF
C3815 _567_/Y _485_/D 2.98fF
C3816 _587_/A _537_/a_227_47# 0.03fF
C3817 _370_/a_68_297# _635_/a_27_413# 0.02fF
C3818 _392_/Y _392_/A 1.55fF
C3819 _390_/B _481_/A 0.19fF
C3820 _510_/A _408_/X 0.01fF
C3821 _607_/X _606_/A 0.01fF
C3822 _374_/a_78_199# VPWR 0.62fF
C3823 output22/a_27_47# M[14] 0.43fF
C3824 _386_/X _446_/X 0.02fF
C3825 B[0] _485_/D 0.03fF
C3826 _386_/a_841_47# _479_/a_68_297# 0.01fF
C3827 _633_/Y _390_/B 0.49fF
C3828 _572_/A _621_/X 0.04fF
C3829 _540_/X _559_/a_539_297# 0.04fF
C3830 _465_/a_109_297# _464_/A 0.01fF
C3831 _616_/B _624_/a_206_369# 0.45fF
C3832 _454_/X _519_/A 0.07fF
C3833 _621_/X _622_/a_29_53# 0.14fF
C3834 _522_/a_76_199# _521_/X 0.22fF
C3835 _378_/A VPWR 2.81fF
C3836 _529_/a_27_47# _531_/C 0.08fF
C3837 _346_/a_161_47# VPWR 1.15fF
C3838 VPWR _537_/a_539_297# 0.02fF
C3839 _484_/a_78_199# _484_/a_292_297# 0.03fF
C3840 VPWR _464_/Y 0.80fF
C3841 _442_/D _483_/a_93_21# 0.04fF
C3842 _557_/a_109_297# VPWR 0.01fF
C3843 _417_/A _367_/C 0.16fF
C3844 _603_/Y _604_/a_209_297# 0.03fF
C3845 _563_/D _530_/X 0.05fF
C3846 _386_/a_62_47# _515_/Y 0.09fF
C3847 B[0] _483_/X 0.15fF
C3848 _458_/X _460_/a_226_47# 0.07fF
C3849 B[1] _328_/A 0.05fF
C3850 _417_/D _514_/A 0.45fF
C3851 B[2] A[2] 0.01fF
C3852 _513_/A _543_/B 0.65fF
C3853 _343_/a_76_199# _343_/a_489_413# 0.12fF
C3854 _560_/a_27_47# _315_/a_161_47# 0.01fF
C3855 _569_/A _595_/a_227_47# 0.30fF
C3856 _428_/a_299_297# VPWR 0.68fF
C3857 _326_/A _411_/A 0.01fF
C3858 A[6] _479_/B 0.09fF
C3859 _419_/a_226_47# VPWR 0.08fF
C3860 _521_/a_292_297# _483_/X 0.02fF
C3861 M[0] _581_/B 0.01fF
C3862 _521_/a_78_199# _488_/X 0.22fF
C3863 _400_/a_80_21# _400_/a_209_297# 0.16fF
C3864 _505_/a_80_21# VPWR 0.33fF
C3865 _583_/a_76_199# _583_/a_489_413# 0.12fF
C3866 _375_/a_448_47# VPWR 0.04fF
C3867 _347_/A _514_/A 0.01fF
C3868 VPWR _316_/a_664_47# 0.37fF
C3869 VPWR _508_/a_539_297# 0.02fF
C3870 _495_/a_226_47# VPWR 0.16fF
C3871 _328_/B _481_/A 0.09fF
C3872 _570_/B _570_/A 0.90fF
C3873 _443_/B VPWR 1.42fF
C3874 _370_/A _370_/B 1.25fF
C3875 _583_/X _607_/a_215_47# 0.08fF
C3876 _371_/A _432_/B 0.08fF
C3877 _513_/A _565_/a_209_297# 0.12fF
C3878 _375_/X _423_/a_215_47# 0.11fF
C3879 _487_/X _381_/B 0.07fF
C3880 _577_/a_226_47# _549_/X 0.02fF
C3881 _378_/a_62_47# _378_/a_558_47# 0.03fF
C3882 _328_/B _633_/Y 0.02fF
C3883 _519_/C _542_/A 0.31fF
C3884 _488_/a_226_47# _559_/a_77_199# 0.00fF
C3885 _538_/Y _486_/X 0.04fF
C3886 _320_/a_161_47# _631_/A 0.68fF
C3887 _521_/X _521_/a_215_47# 0.01fF
C3888 _451_/A _564_/A 0.10fF
C3889 _576_/a_76_199# _530_/X 0.17fF
C3890 _383_/X _332_/a_68_297# 0.14fF
C3891 _362_/a_226_47# _361_/a_76_199# 0.01fF
C3892 _410_/B _446_/X 0.43fF
C3893 _569_/A _627_/C 0.03fF
C3894 _633_/Y _471_/A 0.02fF
C3895 _386_/X _442_/D 1.20fF
C3896 _408_/B _394_/a_381_47# 0.00fF
C3897 _544_/A _516_/A 1.39fF
C3898 _513_/a_27_47# _513_/a_109_47# 0.03fF
C3899 _464_/A _497_/a_68_297# 0.03fF
C3900 _432_/A _430_/A 0.58fF
C3901 _398_/a_226_47# _398_/a_489_413# 0.02fF
C3902 _398_/a_76_199# _398_/a_226_297# 0.01fF
C3903 _542_/B _514_/B 0.42fF
C3904 _365_/a_299_297# VPWR 0.65fF
C3905 _613_/X _442_/D 0.32fF
C3906 _569_/Y B[7] 0.21fF
C3907 _350_/X _398_/X 2.38fF
C3908 _519_/A _337_/A 0.13fF
C3909 B[2] _610_/A 0.52fF
C3910 _542_/A _539_/X 0.05fF
C3911 _328_/A _383_/X 0.40fF
C3912 _614_/a_76_199# _614_/a_226_47# 0.49fF
C3913 _363_/A _343_/X 0.01fF
C3914 _484_/a_215_47# _367_/C 0.11fF
C3915 _381_/C _381_/B 1.99fF
C3916 _608_/X _627_/D 0.21fF
C3917 _526_/a_76_199# _553_/a_78_199# 0.02fF
C3918 _463_/a_76_199# _463_/a_489_413# 0.12fF
C3919 _370_/A _371_/B 0.19fF
C3920 input12/a_381_47# _620_/a_76_199# 0.03fF
C3921 _598_/a_68_297# _598_/B 0.33fF
C3922 _363_/B B[5] 0.25fF
C3923 B[0] _451_/a_27_47# 0.11fF
C3924 _598_/B _599_/Y 0.14fF
C3925 _530_/X _547_/a_222_93# 0.09fF
C3926 _627_/C _627_/D 0.69fF
C3927 _613_/X _588_/Y 0.37fF
C3928 _613_/a_77_199# _433_/Y 0.21fF
C3929 _435_/a_27_47# _566_/Y 0.00fF
C3930 _584_/A _408_/a_68_297# 0.01fF
C3931 _352_/X _631_/A 0.24fF
C3932 _503_/A _588_/A 0.22fF
C3933 _401_/A _558_/X 0.37fF
C3934 _385_/a_381_47# _442_/B 0.18fF
C3935 _567_/B _458_/X 0.24fF
C3936 _359_/a_68_297# _358_/a_27_47# 0.01fF
C3937 _406_/A _631_/B 0.43fF
C3938 _442_/A _469_/X 0.03fF
C3939 _613_/a_77_199# _586_/S 0.27fF
C3940 _417_/A _380_/A 0.03fF
C3941 _381_/B _570_/A 0.67fF
C3942 output26/a_27_47# M[3] 0.47fF
C3943 input3/a_381_47# A[2] 0.02fF
C3944 input3/a_62_47# _390_/D 0.31fF
C3945 _499_/a_299_297# _531_/A 0.03fF
C3946 _566_/A _503_/A 0.03fF
C3947 _494_/a_76_199# _492_/X 0.40fF
C3948 _494_/X VPWR 1.71fF
C3949 _453_/X _485_/D 0.01fF
C3950 output30/a_27_47# _557_/Y 0.22fF
C3951 _557_/Y _558_/a_539_297# 0.02fF
C3952 _542_/C _381_/B 0.09fF
C3953 _623_/a_226_297# _622_/X 0.01fF
C3954 _386_/a_381_47# _386_/a_664_47# 0.09fF
C3955 _458_/X _420_/X 0.01fF
C3956 _410_/B _442_/D 0.05fF
C3957 _535_/Y _472_/B 0.41fF
C3958 _326_/A _409_/a_78_199# 0.13fF
C3959 _584_/a_68_297# _627_/B 0.35fF
C3960 _583_/X input12/a_558_47# 0.15fF
C3961 _544_/A _568_/a_77_199# 0.41fF
C3962 output30/a_27_47# _467_/Y 0.40fF
C3963 _594_/a_109_297# _573_/Y 0.05fF
C3964 _382_/A _542_/D 0.05fF
C3965 _417_/D _449_/A 0.01fF
C3966 _530_/a_489_413# _531_/B 0.19fF
C3967 _608_/a_493_297# _584_/A 0.02fF
C3968 _419_/X _383_/a_76_199# 0.10fF
C3969 _461_/a_78_199# _461_/a_292_297# 0.03fF
C3970 _518_/X _530_/X 0.07fF
C3971 _524_/a_215_47# _525_/a_76_199# 0.01fF
C3972 _367_/C _366_/a_76_199# 0.01fF
C3973 _338_/a_79_199# VPWR 0.65fF
C3974 _487_/X _542_/A 0.18fF
C3975 _587_/A _533_/a_323_297# 0.07fF
C3976 _564_/A _627_/B 0.41fF
C3977 _351_/A VPWR 1.78fF
C3978 _614_/a_76_199# _613_/X 0.32fF
C3979 _614_/a_226_47# _611_/X 0.16fF
C3980 _550_/a_493_297# _521_/X 0.12fF
C3981 _436_/A _510_/A 0.01fF
C3982 _313_/A _442_/B 0.06fF
C3983 _533_/X _510_/X 0.00fF
C3984 _513_/A _454_/X 2.00fF
C3985 _510_/a_68_297# _471_/A 0.01fF
C3986 _510_/a_150_297# _472_/Y 0.01fF
C3987 _410_/a_27_47# _542_/C 0.21fF
C3988 _561_/A _519_/A 0.63fF
C3989 VPWR _621_/a_493_297# 0.01fF
C3990 _381_/B _535_/A 0.45fF
C3991 _513_/A _334_/a_27_47# 0.00fF
C3992 _497_/A _406_/Y 0.02fF
C3993 _580_/B _579_/X 0.19fF
C3994 _563_/A _586_/S 0.02fF
C3995 input12/a_664_47# _620_/X 0.02fF
C3996 input12/a_62_47# _619_/Y 0.01fF
C3997 _627_/X _584_/A 0.11fF
C3998 _590_/A _592_/a_113_297# 0.16fF
C3999 _408_/B _391_/A 0.10fF
C4000 _631_/B _350_/C 0.42fF
C4001 _610_/A _469_/X 1.71fF
C4002 _384_/X _396_/X 1.80fF
C4003 VPWR _397_/a_489_413# 0.45fF
C4004 _358_/a_27_47# _358_/a_109_47# 0.03fF
C4005 _533_/a_227_297# VPWR 0.01fF
C4006 _627_/A _433_/Y 0.67fF
C4007 _544_/A _479_/A 0.03fF
C4008 _519_/a_183_297# _542_/A 0.01fF
C4009 _544_/A _340_/A 1.08fF
C4010 _359_/a_68_297# _359_/B 0.43fF
C4011 _568_/a_77_199# _566_/Y 0.28fF
C4012 _381_/C _542_/A 1.12fF
C4013 _586_/S _627_/A 0.85fF
C4014 _576_/a_556_47# VPWR 0.02fF
C4015 _503_/a_558_47# VPWR 0.22fF
C4016 _569_/Y VPWR 2.45fF
C4017 _547_/X _486_/A 0.54fF
C4018 _506_/Y _533_/a_227_47# 0.07fF
C4019 _363_/A _350_/B 0.08fF
C4020 _544_/A _588_/A 0.66fF
C4021 _631_/B _367_/C 0.48fF
C4022 _360_/a_226_47# _360_/X 0.05fF
C4023 _343_/X _329_/X 1.11fF
C4024 _420_/X _350_/B 0.05fF
C4025 _485_/D _542_/D 0.47fF
C4026 _455_/X _533_/a_77_199# 0.09fF
C4027 _390_/D _547_/X 0.06fF
C4028 _627_/A _540_/X 0.03fF
C4029 _499_/a_81_21# _497_/B 0.02fF
C4030 _544_/A _566_/A 0.45fF
C4031 _543_/B _561_/A 0.00fF
C4032 M[7] _558_/X 0.09fF
C4033 _623_/X _633_/Y 0.05fF
C4034 _448_/A _447_/X 0.23fF
C4035 _533_/X _488_/X 0.29fF
C4036 _519_/X _519_/C 0.01fF
C4037 _542_/A _570_/A 0.03fF
C4038 _533_/a_77_199# _509_/A 0.01fF
C4039 _497_/A _527_/A 0.67fF
C4040 _455_/X _417_/A 0.77fF
C4041 _467_/Y _465_/X 0.66fF
C4042 _461_/a_215_47# _422_/X 0.11fF
C4043 _436_/A _631_/A 0.17fF
C4044 _580_/A _581_/B 0.04fF
C4045 _538_/Y _537_/a_77_199# 0.15fF
C4046 _510_/A _478_/A 0.57fF
C4047 _583_/X _583_/a_76_199# 0.24fF
C4048 _611_/X _613_/X 1.36fF
C4049 _542_/C _542_/A 0.86fF
C4050 _324_/a_841_47# _367_/C 0.05fF
C4051 _490_/a_292_297# VPWR 0.01fF
C4052 _587_/A _475_/a_68_297# 0.37fF
C4053 _540_/X _548_/X 2.39fF
C4054 _599_/A _607_/a_215_47# 0.01fF
C4055 _457_/a_226_47# VPWR 0.10fF
C4056 _411_/B _542_/C 0.13fF
C4057 _347_/A _512_/a_215_47# 0.10fF
C4058 _559_/X _574_/X 0.10fF
C4059 _617_/a_113_297# _616_/Y 0.04fF
C4060 VPWR _500_/a_215_47# 0.07fF
C4061 _576_/X _575_/X 0.38fF
C4062 _559_/X _503_/A 0.04fF
C4063 _335_/a_664_47# VPWR 0.35fF
C4064 output25/a_27_47# _374_/a_78_199# 0.03fF
C4065 _510_/X _509_/Y 0.60fF
C4066 _578_/a_78_199# _559_/X 0.01fF
C4067 _566_/Y _588_/A 0.97fF
C4068 _362_/a_76_199# _362_/a_226_47# 0.49fF
C4069 _509_/Y _511_/a_93_21# 0.56fF
C4070 _448_/A _563_/B 0.06fF
C4071 _534_/a_209_297# _386_/A 0.07fF
C4072 _444_/Y _633_/Y 0.02fF
C4073 _563_/A _378_/A 1.30fF
C4074 input5/a_664_47# _431_/a_226_47# 0.01fF
C4075 input5/a_558_47# _431_/a_489_413# 0.02fF
C4076 input5/a_841_47# _431_/a_76_199# 0.02fF
C4077 _572_/a_68_297# _573_/A 0.27fF
C4078 input2/a_27_47# A[1] 0.40fF
C4079 _567_/Y _570_/X 0.14fF
C4080 _526_/a_226_47# VPWR 0.11fF
C4081 _566_/A _566_/Y 1.73fF
C4082 _460_/a_76_199# VPWR 0.47fF
C4083 _430_/A _371_/A 0.05fF
C4084 _332_/X _366_/a_226_297# 0.03fF
C4085 _542_/A _535_/A 0.03fF
C4086 _603_/Y _555_/a_298_297# 0.15fF
C4087 _426_/a_68_297# _466_/X 0.07fF
C4088 _441_/a_78_199# _340_/A 0.48fF
C4089 _334_/a_27_47# _337_/A 0.18fF
C4090 _351_/a_219_297# _351_/a_27_53# 0.22fF
C4091 _379_/a_493_297# VPWR 0.01fF
C4092 _598_/B _616_/A 1.06fF
C4093 _574_/X _616_/B 1.07fF
C4094 input6/a_27_47# _330_/A 0.07fF
C4095 _625_/a_27_297# _601_/A 0.24fF
C4096 _631_/A _350_/X 0.17fF
C4097 A[6] _542_/D 0.03fF
C4098 _390_/B _558_/X 0.90fF
C4099 _375_/X _382_/B 0.10fF
C4100 _423_/X _390_/B 0.54fF
C4101 _347_/A _417_/D 2.15fF
C4102 _518_/a_256_47# _381_/B 0.04fF
C4103 _383_/X _397_/a_226_47# 0.01fF
C4104 _520_/a_489_413# VPWR 0.39fF
C4105 _382_/X _383_/X 0.01fF
C4106 _347_/a_27_47# _380_/A 0.01fF
C4107 _549_/a_76_199# _559_/X 0.07fF
C4108 _478_/A _483_/X 0.01fF
C4109 _519_/A VPWR 7.23fF
C4110 _442_/a_27_47# _442_/a_109_47# 0.03fF
C4111 _417_/A _452_/A 0.53fF
C4112 _406_/A _458_/a_292_297# 0.02fF
C4113 _542_/a_27_47# _542_/a_109_47# 0.03fF
C4114 _584_/a_68_297# VPWR 0.29fF
C4115 _616_/Y _601_/A 0.58fF
C4116 _591_/Y _588_/A 0.43fF
C4117 _348_/a_27_47# _328_/A 0.07fF
C4118 _602_/Y _604_/a_80_21# 0.24fF
C4119 _353_/X _359_/B 0.02fF
C4120 _380_/A _631_/B 0.11fF
C4121 _611_/a_27_297# B[7] 0.26fF
C4122 _615_/a_78_199# VPWR 0.80fF
C4123 _353_/X _353_/a_68_297# 0.27fF
C4124 _455_/X _469_/X 0.03fF
C4125 B[1] _335_/a_558_47# 0.20fF
C4126 _375_/X _330_/A 0.32fF
C4127 _443_/B _470_/a_80_21# 0.30fF
C4128 input12/a_664_47# VPWR 0.35fF
C4129 _465_/X _427_/A 0.05fF
C4130 _586_/a_439_47# _622_/C 0.03fF
C4131 _517_/X _515_/A 0.18fF
C4132 _511_/X _550_/a_78_199# 0.33fF
C4133 _324_/a_381_47# _324_/a_558_47# 0.32fF
C4134 _541_/a_493_297# VPWR 0.02fF
C4135 _564_/A VPWR 1.80fF
C4136 _509_/A _469_/X 0.34fF
C4137 _408_/a_68_297# _408_/a_150_297# 0.02fF
C4138 _533_/X _511_/X 0.24fF
C4139 _445_/A _409_/a_78_199# 0.30fF
C4140 _356_/a_78_199# _481_/A 0.25fF
C4141 _422_/a_226_297# _412_/X 0.01fF
C4142 _567_/B _587_/A 0.27fF
C4143 _549_/X _575_/X 0.01fF
C4144 _387_/a_493_297# _633_/Y 0.02fF
C4145 _487_/X _488_/a_489_413# 0.22fF
C4146 _513_/A _561_/A 0.05fF
C4147 _506_/A _442_/D 0.03fF
C4148 _418_/a_68_297# _418_/B 0.30fF
C4149 _424_/a_489_413# _422_/X 0.11fF
C4150 _353_/a_68_297# _353_/a_150_297# 0.02fF
C4151 _578_/a_78_199# _550_/X 0.13fF
C4152 _374_/a_78_199# _374_/a_292_297# 0.03fF
C4153 _473_/a_77_199# _473_/a_227_47# 0.24fF
C4154 _502_/a_78_199# _468_/X 0.49fF
C4155 VPWR _507_/Y 2.72fF
C4156 _519_/A _314_/X 0.03fF
C4157 _480_/Y _482_/X 0.91fF
C4158 _318_/a_303_47# _485_/A 0.03fF
C4159 _573_/A _588_/A 0.25fF
C4160 _536_/Y _487_/X 0.02fF
C4161 _557_/Y _530_/X 0.22fF
C4162 _369_/a_76_199# _343_/X 0.22fF
C4163 _543_/B VPWR 4.64fF
C4164 _602_/A _530_/X 0.53fF
C4165 _411_/a_68_297# _470_/a_209_297# 0.00fF
C4166 _363_/A _371_/B 0.16fF
C4167 _519_/X _381_/C 1.23fF
C4168 _456_/a_76_199# _456_/a_226_47# 0.49fF
C4169 _561_/A _454_/X 0.03fF
C4170 _451_/A _627_/B 0.16fF
C4171 _543_/B _544_/a_664_47# 0.08fF
C4172 _543_/Y _544_/a_381_47# 0.01fF
C4173 _587_/A _468_/a_78_199# 0.26fF
C4174 input9/a_27_47# VPWR 0.53fF
C4175 _568_/a_227_47# _570_/B 0.04fF
C4176 _396_/a_584_47# _330_/A 0.02fF
C4177 _628_/Y output23/a_27_47# 0.41fF
C4178 _412_/X _421_/X 2.44fF
C4179 _467_/Y _530_/X 0.03fF
C4180 _442_/a_27_47# _316_/a_841_47# 0.01fF
C4181 _565_/a_209_297# VPWR 0.46fF
C4182 _500_/a_292_297# VPWR 0.05fF
C4183 B[7] _454_/X 0.71fF
C4184 _543_/A _514_/a_68_297# 0.20fF
C4185 _350_/X _391_/a_68_297# 0.20fF
C4186 _628_/a_382_297# _628_/a_28_47# 0.03fF
C4187 _516_/A _482_/X 0.06fF
C4188 _476_/a_250_297# _390_/B 0.17fF
C4189 _482_/X _539_/A 0.06fF
C4190 _408_/B _442_/B 1.33fF
C4191 _469_/A _545_/Y 0.20fF
C4192 _545_/Y _544_/a_841_47# 0.01fF
C4193 _418_/B _542_/D 1.87fF
C4194 _584_/A _394_/a_62_47# 0.38fF
C4195 _566_/Y _559_/X 0.03fF
C4196 _557_/A _401_/A 0.37fF
C4197 _595_/X _593_/Y 0.71fF
C4198 _538_/Y VPWR 1.53fF
C4199 _443_/A _346_/A 0.09fF
C4200 _423_/a_78_199# _631_/A 0.18fF
C4201 _561_/A _451_/A 0.05fF
C4202 _455_/a_79_199# _378_/A 0.01fF
C4203 _488_/a_489_413# _570_/A 0.00fF
C4204 _379_/a_78_199# _417_/A 0.18fF
C4205 _327_/a_215_47# _328_/B 0.17fF
C4206 _569_/A _469_/X 0.78fF
C4207 _382_/A _383_/a_76_199# 0.01fF
C4208 _451_/A B[7] 0.15fF
C4209 _626_/Y _522_/a_226_297# 0.02fF
C4210 _433_/a_397_297# VPWR 0.57fF
C4211 _497_/B _497_/A 0.40fF
C4212 _613_/a_227_47# _586_/a_505_21# 0.03fF
C4213 _509_/Y _511_/X 0.38fF
C4214 _583_/a_226_47# VPWR 0.09fF
C4215 _628_/a_382_297# _622_/X 0.00fF
C4216 _583_/X _581_/a_27_93# 0.06fF
C4217 _365_/a_81_21# _629_/X 0.01fF
C4218 _536_/Y _570_/A 0.40fF
C4219 _442_/D _515_/A 0.12fF
C4220 _473_/a_227_47# _471_/A 0.05fF
C4221 _503_/A _530_/X 0.03fF
C4222 _574_/X _530_/X 1.13fF
C4223 _419_/a_76_199# _419_/a_226_297# 0.01fF
C4224 _419_/a_226_47# _419_/a_489_413# 0.02fF
C4225 _455_/a_222_93# _419_/a_76_199# 0.00fF
C4226 _455_/a_79_199# _419_/a_226_47# 0.00fF
C4227 _570_/B _485_/D 0.71fF
C4228 _578_/a_78_199# _530_/X 0.11fF
C4229 A[5] _630_/X 0.82fF
C4230 _611_/a_27_297# VPWR 0.64fF
C4231 _627_/a_27_297# _627_/a_109_297# 0.02fF
C4232 _626_/Y _485_/D 0.03fF
C4233 _410_/a_197_47# _410_/C 0.09fF
C4234 _505_/a_80_21# _505_/a_209_297# 0.16fF
C4235 _540_/a_250_297# _469_/X 0.10fF
C4236 _613_/a_323_297# _627_/D 0.12fF
C4237 _557_/Y _557_/B 0.94fF
C4238 _542_/D _627_/a_277_297# 0.01fF
C4239 _566_/A _571_/a_256_47# 0.03fF
C4240 _500_/a_215_47# _531_/C 0.01fF
C4241 _573_/Y _585_/B 0.06fF
C4242 _469_/a_62_47# _586_/a_76_199# 0.00fF
C4243 _566_/Y _571_/a_93_21# 0.01fF
C4244 _585_/B _544_/a_381_47# 0.00fF
C4245 _468_/a_215_47# _390_/B 0.11fF
C4246 _351_/X _363_/B 0.03fF
C4247 _375_/X _442_/B 1.63fF
C4248 _311_/a_27_47# _449_/A 0.04fF
C4249 _538_/Y _559_/a_539_297# 0.03fF
C4250 _316_/a_664_47# _316_/a_841_47# 0.29fF
C4251 _527_/B _527_/A 1.61fF
C4252 _583_/X _622_/C 0.01fF
C4253 _467_/Y _557_/B 0.74fF
C4254 _495_/a_76_199# _495_/a_226_297# 0.01fF
C4255 _495_/a_226_47# _495_/a_489_413# 0.02fF
C4256 VPWR _486_/X 4.97fF
C4257 _510_/A _385_/a_62_47# 0.14fF
C4258 _476_/X _492_/X 0.03fF
C4259 _539_/A _539_/X 0.56fF
C4260 _412_/a_76_199# _437_/a_79_199# 0.04fF
C4261 _595_/a_77_199# _595_/a_227_47# 0.24fF
C4262 _386_/a_558_47# VPWR 0.24fF
C4263 _622_/C _622_/X 0.01fF
C4264 _628_/a_734_297# B[7] 0.13fF
C4265 M[14] _466_/X 0.00fF
C4266 _491_/a_489_413# VPWR 0.39fF
C4267 _536_/Y _535_/A 0.24fF
C4268 _513_/A VPWR 8.66fF
C4269 _581_/a_27_93# _580_/a_68_297# 0.00fF
C4270 _408_/X _394_/a_664_47# 0.02fF
C4271 _543_/Y _546_/a_226_297# 0.02fF
C4272 _566_/A _546_/a_226_47# 0.06fF
C4273 B[1] _326_/A 0.43fF
C4274 _361_/a_489_413# _374_/X 0.13fF
C4275 _569_/Y _627_/A 0.14fF
C4276 _503_/a_558_47# _627_/A 0.11fF
C4277 _351_/A _351_/a_27_53# 0.18fF
C4278 _390_/D _481_/A 0.50fF
C4279 _597_/a_493_297# VPWR 0.01fF
C4280 _347_/A _477_/a_78_199# 0.28fF
C4281 _591_/Y _616_/B 0.03fF
C4282 _519_/A _484_/a_292_297# 0.07fF
C4283 _534_/a_80_21# _534_/a_303_47# 0.04fF
C4284 _425_/a_76_199# _424_/X 0.24fF
C4285 _390_/D _633_/Y 0.07fF
C4286 _612_/Y _633_/Y 0.03fF
C4287 _556_/Y _557_/Y 1.45fF
C4288 _552_/a_76_199# _554_/A 0.24fF
C4289 _472_/Y _478_/A 0.80fF
C4290 _452_/A _631_/B 0.00fF
C4291 _454_/X VPWR 10.26fF
C4292 _334_/a_27_47# VPWR 0.80fF
C4293 _544_/A _448_/B 2.82fF
C4294 _510_/X _533_/a_77_199# 0.38fF
C4295 _563_/D _408_/B 0.70fF
C4296 _417_/D _518_/a_93_21# 0.10fF
C4297 _487_/X _480_/Y 0.12fF
C4298 _479_/A _482_/X 0.13fF
C4299 _533_/a_77_199# _511_/a_93_21# 0.04fF
C4300 _381_/B _485_/D 1.30fF
C4301 _556_/Y _467_/Y 0.00fF
C4302 _557_/A M[7] 0.34fF
C4303 B[7] _627_/B 0.88fF
C4304 _436_/A _437_/X 0.00fF
C4305 _419_/X _420_/a_222_93# 0.13fF
C4306 _336_/a_78_199# _332_/X 0.18fF
C4307 _365_/a_81_21# _432_/B 0.19fF
C4308 _455_/a_448_47# _413_/X 0.17fF
C4309 _469_/a_558_47# _584_/A 0.10fF
C4310 _347_/A _518_/a_93_21# 0.05fF
C4311 _386_/A _385_/a_558_47# 0.11fF
C4312 _544_/A _530_/X 0.25fF
C4313 _553_/a_493_297# _525_/X 0.02fF
C4314 _393_/A _363_/A 1.02fF
C4315 _563_/a_27_297# _563_/a_277_297# 0.05fF
C4316 _485_/a_197_47# _542_/D 0.07fF
C4317 _553_/a_215_47# _504_/X 0.03fF
C4318 _494_/a_76_199# _626_/Y 0.08fF
C4319 _631_/B _421_/X 0.17fF
C4320 _329_/a_226_47# _328_/X 0.53fF
C4321 _393_/A _420_/X 0.11fF
C4322 _384_/X _423_/X 0.03fF
C4323 _590_/B _572_/A 0.13fF
C4324 _504_/a_227_47# _390_/B 0.11fF
C4325 _458_/X _439_/a_556_47# 0.02fF
C4326 _328_/A _481_/A 0.03fF
C4327 _451_/A VPWR 2.62fF
C4328 _495_/a_226_297# _468_/X 0.01fF
C4329 _495_/a_489_413# _494_/X 0.14fF
C4330 _584_/A _449_/A 0.01fF
C4331 _516_/A _487_/X 1.13fF
C4332 _426_/A _371_/B 0.39fF
C4333 _563_/D _445_/a_68_297# 0.43fF
C4334 _381_/B _483_/X 0.03fF
C4335 _487_/X _539_/A 3.19fF
C4336 B[1] _633_/a_265_297# 0.03fF
C4337 _633_/Y _328_/A 0.03fF
C4338 _561_/A B[7] 0.03fF
C4339 _383_/X _447_/B 0.10fF
C4340 _436_/A _439_/a_76_199# 0.00fF
C4341 _447_/a_68_297# _417_/a_27_47# 0.01fF
C4342 _356_/a_215_47# _447_/B 0.08fF
C4343 _408_/B _336_/a_292_297# 0.08fF
C4344 _476_/a_250_297# _504_/a_77_199# 0.08fF
C4345 _393_/A _411_/A 0.08fF
C4346 _591_/Y _592_/a_113_297# 0.04fF
C4347 _360_/X B[5] 0.03fF
C4348 _543_/Y _469_/a_841_47# 0.00fF
C4349 _573_/Y _572_/B 0.05fF
C4350 _530_/X _504_/X 0.08fF
C4351 _431_/a_226_47# _431_/a_489_413# 0.02fF
C4352 _431_/a_76_199# _431_/a_226_297# 0.01fF
C4353 _327_/a_292_297# VPWR 0.01fF
C4354 _461_/a_215_47# _406_/Y 0.27fF
C4355 _634_/Y _635_/Y 0.09fF
C4356 _516_/A _381_/C 0.58fF
C4357 _341_/a_27_47# VPWR 0.66fF
C4358 _469_/A _522_/X 0.01fF
C4359 _527_/a_109_297# VPWR 0.01fF
C4360 _585_/B _403_/a_27_47# 0.29fF
C4361 _338_/X _337_/X 0.00fF
C4362 _417_/A _475_/A 0.03fF
C4363 _566_/Y _530_/X 0.50fF
C4364 _482_/a_68_297# _477_/a_215_47# 0.02fF
C4365 _473_/a_323_297# VPWR 0.02fF
C4366 _517_/a_68_297# _520_/X 0.01fF
C4367 _476_/a_93_21# _587_/A 0.05fF
C4368 _337_/A VPWR 6.94fF
C4369 _542_/C _480_/Y 0.09fF
C4370 _369_/a_76_199# _370_/B 0.24fF
C4371 _556_/Y _606_/A 0.04fF
C4372 _613_/a_227_47# _590_/A 0.02fF
C4373 _400_/a_80_21# _420_/X 0.10fF
C4374 _411_/B _437_/a_222_93# 0.30fF
C4375 _329_/a_226_47# _329_/X 0.05fF
C4376 A[6] _381_/B 1.11fF
C4377 _361_/a_76_199# _374_/X 0.18fF
C4378 _628_/a_734_297# VPWR 0.45fF
C4379 _417_/D _311_/a_27_47# 0.00fF
C4380 _442_/D A[3] 0.03fF
C4381 _630_/X _398_/X 0.75fF
C4382 B[2] _597_/a_78_199# 0.05fF
C4383 _581_/a_206_47# VPWR 0.00fF
C4384 _411_/B _510_/A 0.31fF
C4385 _417_/D _410_/C 0.03fF
C4386 _538_/A _469_/X 1.15fF
C4387 _628_/a_300_47# _623_/X 0.12fF
C4388 _628_/a_28_47# _625_/Y 0.17fF
C4389 _510_/X _469_/X 1.00fF
C4390 _583_/X _612_/A 0.05fF
C4391 _370_/A _635_/a_384_47# 0.13fF
C4392 _516_/A _570_/A 2.23fF
C4393 _589_/a_76_199# _589_/a_489_413# 0.12fF
C4394 _511_/a_93_21# _469_/X 0.31fF
C4395 _586_/S _541_/a_215_47# 0.01fF
C4396 _349_/a_78_199# _351_/A 0.23fF
C4397 _358_/a_303_47# _381_/B 0.05fF
C4398 _408_/a_68_297# _394_/a_381_47# 0.02fF
C4399 _347_/A _410_/C 0.15fF
C4400 _516_/A _542_/C 0.17fF
C4401 _504_/a_77_199# _468_/a_215_47# 0.02fF
C4402 _539_/A _508_/a_77_199# 0.44fF
C4403 _465_/a_27_297# _465_/X 0.21fF
C4404 _386_/X _392_/A 0.69fF
C4405 _542_/C _539_/A 0.03fF
C4406 _417_/a_197_47# _447_/X 0.03fF
C4407 _571_/a_93_21# _571_/a_256_47# 0.03fF
C4408 _542_/A _485_/D 1.56fF
C4409 _453_/a_584_47# _542_/D 0.02fF
C4410 _588_/Y A[3] 0.06fF
C4411 _543_/A _433_/Y 0.04fF
C4412 input3/a_558_47# _485_/D 0.07fF
C4413 _627_/A _507_/Y 0.09fF
C4414 _478_/a_27_47# _505_/a_80_21# 0.01fF
C4415 _381_/a_27_47# _358_/a_27_47# 0.02fF
C4416 _567_/B _433_/Y 0.50fF
C4417 _466_/X _467_/a_481_47# 0.06fF
C4418 _543_/B _627_/A 0.39fF
C4419 _595_/a_323_297# VPWR 0.02fF
C4420 VPWR _627_/B 9.70fF
C4421 _537_/a_77_199# VPWR 0.91fF
C4422 _625_/Y _622_/X 0.04fF
C4423 _583_/X _601_/Y 0.18fF
C4424 _542_/A _483_/X 0.72fF
C4425 _320_/a_161_47# _367_/C 0.00fF
C4426 _539_/A _535_/A 0.01fF
C4427 input4/a_27_47# _483_/X 0.10fF
C4428 _382_/a_68_297# _452_/A 0.07fF
C4429 _620_/X VPWR 2.51fF
C4430 _433_/a_109_47# _629_/B 0.00fF
C4431 _475_/X _587_/A 0.65fF
C4432 _487_/X _479_/A 0.31fF
C4433 _487_/X _340_/A 0.16fF
C4434 _455_/X _533_/a_227_47# 0.19fF
C4435 _363_/B _398_/X 0.20fF
C4436 _567_/B _540_/X 0.58fF
C4437 _506_/Y _478_/A 0.10fF
C4438 _452_/a_68_297# _452_/A 0.35fF
C4439 _513_/a_303_47# _542_/A 0.03fF
C4440 _476_/X _456_/X 0.03fF
C4441 _533_/a_77_199# _511_/X 0.02fF
C4442 _411_/a_68_297# _633_/Y 0.01fF
C4443 _524_/a_78_199# _524_/X 0.22fF
C4444 _561_/A VPWR 6.66fF
C4445 B[1] _445_/A 0.65fF
C4446 _417_/D _584_/A 1.30fF
C4447 _538_/Y _627_/A 0.03fF
C4448 _610_/A _599_/Y 0.06fF
C4449 _347_/A _445_/X 0.16fF
C4450 _634_/Y _370_/B 0.27fF
C4451 B[7] VPWR 12.03fF
C4452 _516_/A _413_/X 0.02fF
C4453 _568_/a_77_199# _570_/A 0.01fF
C4454 _589_/a_489_413# _612_/A 0.07fF
C4455 _338_/a_79_199# _338_/a_222_93# 0.51fF
C4456 _544_/A _514_/B 0.52fF
C4457 _347_/A _584_/A 0.13fF
C4458 _422_/X _406_/A 0.16fF
C4459 _545_/Y _547_/X 0.01fF
C4460 _483_/a_256_47# _542_/A 0.01fF
C4461 _476_/X _478_/A 0.19fF
C4462 _477_/a_78_199# _518_/a_93_21# 0.01fF
C4463 B[1] _350_/B 0.90fF
C4464 _429_/a_226_47# _371_/B 0.02fF
C4465 _381_/C _340_/A 0.01fF
C4466 B[2] _601_/A 0.03fF
C4467 _469_/a_381_47# _503_/A 0.06fF
C4468 _410_/C _445_/a_150_297# 0.02fF
C4469 A[6] _542_/A 3.74fF
C4470 _504_/a_77_199# _504_/a_227_47# 0.24fF
C4471 _589_/a_226_47# VPWR 0.10fF
C4472 A[6] input4/a_27_47# 0.09fF
C4473 _526_/a_226_47# _523_/X 0.00fF
C4474 _376_/X _383_/a_489_413# 0.06fF
C4475 _430_/A _363_/a_68_297# 0.27fF
C4476 _381_/a_27_47# _359_/B 0.01fF
C4477 _369_/a_226_297# B[5] 0.01fF
C4478 _534_/a_209_297# _515_/A 0.15fF
C4479 _432_/X _466_/X 0.01fF
C4480 _396_/X _397_/a_226_47# 0.56fF
C4481 _429_/a_76_199# VPWR 0.49fF
C4482 _612_/Y _585_/B 0.16fF
C4483 _623_/X _589_/a_226_297# 0.01fF
C4484 _487_/X _521_/a_493_297# 0.08fF
C4485 _390_/D _585_/B 0.10fF
C4486 VPWR _574_/a_81_21# 0.43fF
C4487 _458_/a_292_297# _421_/X 0.08fF
C4488 _570_/B _570_/X 0.01fF
C4489 _631_/A _366_/a_226_47# 0.01fF
C4490 _459_/a_76_199# _458_/X 0.28fF
C4491 _445_/A _383_/X 0.03fF
C4492 _340_/A _570_/A 0.05fF
C4493 _513_/A _563_/A 1.03fF
C4494 _634_/Y _371_/B 0.67fF
C4495 _596_/a_489_413# _594_/X 0.18fF
C4496 _596_/a_226_47# _595_/X 0.51fF
C4497 _442_/D _442_/B 0.11fF
C4498 _542_/B _442_/D 0.07fF
C4499 _627_/A _486_/X 0.03fF
C4500 _563_/D _517_/X 0.05fF
C4501 _436_/A _406_/A 0.14fF
C4502 _633_/Y _631_/Y 0.07fF
C4503 _410_/a_197_47# _410_/B 0.03fF
C4504 _386_/A _417_/D 0.38fF
C4505 _559_/X _539_/X 0.00fF
C4506 _386_/X _392_/Y 0.66fF
C4507 _425_/a_76_199# _425_/a_489_413# 0.12fF
C4508 _383_/X _350_/B 0.03fF
C4509 _598_/B _593_/A 0.61fF
C4510 _520_/X _472_/B 0.22fF
C4511 _596_/a_76_199# _596_/a_489_413# 0.12fF
C4512 _504_/a_323_297# VPWR 0.02fF
C4513 _347_/A _386_/A 0.16fF
C4514 _516_/A _477_/a_493_297# 0.01fF
C4515 _487_/a_215_47# _454_/X 0.01fF
C4516 _487_/a_78_199# _453_/X 0.30fF
C4517 _566_/A _570_/A 0.03fF
C4518 _563_/A _454_/X 0.03fF
C4519 _350_/C _409_/a_493_297# 0.06fF
C4520 _503_/a_381_47# _503_/a_841_47# 0.03fF
C4521 _503_/a_558_47# _503_/a_664_47# 0.60fF
C4522 _508_/a_227_47# _507_/Y 0.05fF
C4523 _563_/A _334_/a_27_47# 0.22fF
C4524 _631_/B _475_/A 1.24fF
C4525 _392_/A _395_/X 0.30fF
C4526 _417_/D _521_/X 0.15fF
C4527 _511_/X _469_/X 0.02fF
C4528 _538_/Y _537_/a_227_47# 0.02fF
C4529 _579_/a_59_75# M[0] 0.14fF
C4530 _350_/X _399_/a_78_199# 0.33fF
C4531 _566_/A _542_/C 0.08fF
C4532 input10/a_27_47# _429_/a_489_413# 0.02fF
C4533 _390_/B _531_/A 0.00fF
C4534 _481_/a_27_47# _481_/A 0.32fF
C4535 _425_/a_226_47# VPWR 0.15fF
C4536 _440_/a_226_47# _478_/A 0.14fF
C4537 _627_/A _454_/X 0.03fF
C4538 _578_/a_215_47# _551_/a_76_199# 0.01fF
C4539 _439_/X _436_/A 0.01fF
C4540 VPWR _501_/a_109_47# 0.25fF
C4541 _373_/Y VPWR 0.81fF
C4542 output31/a_27_47# M[8] 0.43fF
C4543 _469_/A _587_/A 0.25fF
C4544 _519_/X _485_/D 0.27fF
C4545 _390_/B _469_/X 0.57fF
C4546 _453_/a_93_21# _453_/a_346_47# 0.05fF
C4547 _469_/A _612_/A 0.05fF
C4548 output24/a_27_47# _633_/Y 0.63fF
C4549 _547_/X _486_/a_68_297# 0.01fF
C4550 _570_/X _381_/B 0.28fF
C4551 _475_/A _411_/X 0.12fF
C4552 _563_/B _486_/A 0.01fF
C4553 _605_/a_80_21# _556_/Y 0.15fF
C4554 _631_/A _337_/X 0.02fF
C4555 M[5] _350_/X 0.06fF
C4556 _418_/B _542_/A 0.04fF
C4557 _629_/A _629_/a_68_297# 0.35fF
C4558 _518_/a_250_297# _517_/X 0.10fF
C4559 _612_/Y _616_/Y 0.88fF
C4560 _436_/A _350_/C 0.58fF
C4561 _513_/a_27_47# _542_/B 0.29fF
C4562 _566_/A _535_/A 0.14fF
C4563 _380_/A _352_/X 0.04fF
C4564 _536_/Y _485_/D 0.30fF
C4565 _410_/a_27_47# _446_/a_250_297# 0.02fF
C4566 M[8] _501_/a_481_47# 0.01fF
C4567 _544_/a_664_47# VPWR 0.35fF
C4568 _594_/a_27_297# _615_/a_78_199# 0.01fF
C4569 _524_/a_78_199# _491_/X 0.23fF
C4570 _487_/X _559_/X 0.00fF
C4571 _544_/a_558_47# _544_/a_841_47# 0.07fF
C4572 _633_/Y _490_/a_78_199# 0.13fF
C4573 _630_/X _398_/a_556_47# 0.02fF
C4574 _365_/a_299_297# _363_/A 0.12fF
C4575 _488_/a_226_47# _488_/X 0.05fF
C4576 _606_/Y VPWR 2.59fF
C4577 VPWR _514_/a_150_297# 0.00fF
C4578 _443_/B _411_/A 0.04fF
C4579 input2/a_27_47# _558_/X 0.14fF
C4580 _335_/a_558_47# _633_/Y 0.08fF
C4581 _375_/X _384_/a_489_413# 0.07fF
C4582 _544_/A _378_/a_62_47# 0.41fF
C4583 _374_/a_78_199# _374_/X 0.33fF
C4584 _386_/X _417_/D 0.08fF
C4585 _503_/a_558_47# _475_/a_68_297# 0.01fF
C4586 _478_/A _428_/X 0.36fF
C4587 input14/a_27_47# B[5] 0.45fF
C4588 _431_/a_76_199# _430_/X 0.29fF
C4589 _613_/a_77_199# _627_/B 0.01fF
C4590 _501_/a_109_47# _501_/Y 0.47fF
C4591 B[1] _371_/B 0.10fF
C4592 M[8] _626_/Y 0.03fF
C4593 _386_/X _347_/A 0.24fF
C4594 output31/a_27_47# _465_/a_109_297# 0.03fF
C4595 _567_/B _494_/X 0.34fF
C4596 _585_/B _508_/a_323_297# 0.10fF
C4597 _496_/a_215_47# VPWR 0.07fF
C4598 _314_/X VPWR 1.03fF
C4599 _577_/a_76_199# _577_/a_489_413# 0.12fF
C4600 _601_/Y _599_/A 0.03fF
C4601 _542_/D _367_/C 0.07fF
C4602 _579_/X output17/a_27_47# 0.01fF
C4603 _390_/B _470_/a_209_47# 0.05fF
C4604 B[1] _326_/a_27_47# 0.10fF
C4605 _439_/X _478_/A 0.03fF
C4606 _627_/A _473_/a_323_297# 0.04fF
C4607 _490_/a_78_199# _490_/a_215_47# 0.26fF
C4608 VPWR _559_/a_539_297# 0.02fF
C4609 _476_/X _626_/Y 0.21fF
C4610 input3/a_62_47# _618_/Y 0.01fF
C4611 _548_/a_226_47# _485_/D 0.16fF
C4612 _471_/A _469_/X 0.10fF
C4613 _457_/a_76_199# _457_/a_226_297# 0.01fF
C4614 _457_/a_226_47# _457_/a_489_413# 0.02fF
C4615 VPWR _501_/Y 5.13fF
C4616 _561_/a_27_47# _542_/A 0.23fF
C4617 _610_/A _616_/A 0.51fF
C4618 _469_/A _559_/a_323_297# 0.04fF
C4619 _350_/C _350_/X 0.12fF
C4620 _519_/X A[6] 1.44fF
C4621 _335_/a_664_47# _335_/a_841_47# 0.29fF
C4622 _554_/X _554_/a_68_297# 0.35fF
C4623 _517_/X _518_/X 0.07fF
C4624 _340_/A _477_/a_493_297# 0.04fF
C4625 _329_/a_489_413# VPWR 0.33fF
C4626 _613_/a_77_199# B[7] 0.17fF
C4627 _610_/A _572_/A 0.15fF
C4628 _411_/B _446_/a_250_297# 0.09fF
C4629 _525_/a_226_47# _492_/a_76_199# 0.01fF
C4630 _525_/a_76_199# _492_/a_226_47# 0.01fF
C4631 _559_/X _570_/A 0.01fF
C4632 _563_/A _627_/B 0.25fF
C4633 _547_/X _486_/B 0.26fF
C4634 _583_/X _433_/Y 0.01fF
C4635 _482_/a_150_297# A[6] 0.02fF
C4636 _392_/Y _395_/X 0.03fF
C4637 _394_/a_62_47# _394_/a_381_47# 0.08fF
C4638 _460_/X _462_/a_76_199# 0.46fF
C4639 _496_/a_78_199# _406_/Y 0.48fF
C4640 _342_/X VPWR 3.02fF
C4641 _351_/A _363_/A 0.03fF
C4642 _433_/Y _622_/X 0.77fF
C4643 _526_/a_76_199# _526_/a_226_297# 0.01fF
C4644 _526_/a_226_47# _526_/a_489_413# 0.02fF
C4645 _460_/a_76_199# _460_/a_226_47# 0.49fF
C4646 _360_/X _351_/X 0.17fF
C4647 _351_/A _420_/X 0.03fF
C4648 _326_/a_27_47# _383_/X 0.12fF
C4649 VPWR _466_/a_292_297# 0.01fF
C4650 _627_/A _595_/a_323_297# 0.09fF
C4651 _627_/A _627_/B 0.24fF
C4652 _337_/A _368_/A 0.06fF
C4653 _442_/A _346_/A 0.58fF
C4654 _523_/a_76_199# _511_/X 0.44fF
C4655 _410_/B _347_/A 0.13fF
C4656 _568_/a_227_47# _435_/a_27_47# 0.04fF
C4657 _390_/D _537_/a_323_297# 0.03fF
C4658 _569_/Y _567_/B 0.02fF
C4659 _478_/A _442_/A 0.26fF
C4660 _569_/A _567_/Y 0.02fF
C4661 _563_/A _561_/A 0.28fF
C4662 _329_/a_489_413# _314_/X 0.07fF
C4663 _610_/A _542_/D 0.01fF
C4664 _356_/a_493_297# VPWR 0.01fF
C4665 _442_/D _591_/A 0.12fF
C4666 _426_/A _464_/Y 0.06fF
C4667 _516_/A _382_/A 0.01fF
C4668 _514_/A _515_/A 0.03fF
C4669 _454_/a_76_199# _628_/Y 0.17fF
C4670 _503_/A _472_/B 0.35fF
C4671 _571_/a_93_21# _570_/A 0.00fF
C4672 _436_/A _380_/A 1.18fF
C4673 _627_/D _599_/Y 0.53fF
C4674 _515_/Y _518_/a_584_47# 0.01fF
C4675 _633_/A _632_/a_78_199# 0.23fF
C4676 VPWR _399_/a_215_47# 0.04fF
C4677 _452_/A _320_/a_161_47# 0.58fF
C4678 _627_/C _612_/Y 0.66fF
C4679 _411_/B _437_/X 0.02fF
C4680 _564_/a_219_297# _564_/a_301_297# 0.02fF
C4681 _425_/a_76_199# _407_/Y 0.38fF
C4682 _342_/X _314_/X 0.18fF
C4683 _530_/X _556_/A 0.48fF
C4684 _385_/a_381_47# _394_/a_558_47# 0.04fF
C4685 _440_/X _493_/a_215_47# 0.03fF
C4686 _510_/X _533_/a_227_47# 0.14fF
C4687 _328_/B _631_/B 0.80fF
C4688 _475_/X _433_/Y 0.03fF
C4689 _428_/a_299_297# _426_/A 0.12fF
C4690 _380_/A _542_/D 0.00fF
C4691 _504_/a_77_199# _469_/X 0.01fF
C4692 _368_/B _634_/a_300_297# 0.22fF
C4693 _532_/a_76_199# _532_/a_489_47# 0.14fF
C4694 _588_/Y _591_/A 0.39fF
C4695 _627_/A B[7] 0.04fF
C4696 _520_/X _517_/X 0.49fF
C4697 _360_/X A[5] 0.01fF
C4698 _590_/B _593_/A 0.01fF
C4699 _436_/A _384_/a_226_47# 0.08fF
C4700 _580_/A _579_/a_59_75# 0.25fF
C4701 _527_/B _532_/a_76_199# 0.25fF
C4702 _501_/a_109_47# _531_/C 0.56fF
C4703 _445_/X _410_/C 0.39fF
C4704 _360_/X _419_/X 0.03fF
C4705 _563_/a_27_297# _563_/B 0.41fF
C4706 _584_/a_68_297# _584_/a_150_297# 0.02fF
C4707 input10/a_27_47# _417_/A 0.22fF
C4708 _584_/A _410_/C 0.03fF
C4709 B[7] _548_/X 0.00fF
C4710 _519_/C _453_/a_93_21# 0.29fF
C4711 _326_/A _481_/A 0.63fF
C4712 _615_/a_78_199# _615_/a_292_297# 0.03fF
C4713 VPWR _484_/a_292_297# 0.01fF
C4714 _633_/Y _326_/A 0.18fF
C4715 _516_/A _485_/D 0.27fF
C4716 VPWR _531_/C 4.19fF
C4717 _480_/Y _483_/X 0.02fF
C4718 _481_/A _447_/B 0.19fF
C4719 _487_/X _530_/X 0.05fF
C4720 _574_/X _548_/a_489_413# 0.01fF
C4721 _549_/X _552_/a_76_199# 0.02fF
C4722 _550_/X _552_/a_226_47# 0.00fF
C4723 _329_/a_76_199# _417_/A 0.05fF
C4724 _551_/X _552_/a_489_413# 0.17fF
C4725 _533_/X _552_/a_226_297# 0.03fF
C4726 _613_/a_77_199# VPWR 0.95fF
C4727 _400_/a_209_297# VPWR 0.42fF
C4728 _335_/a_664_47# _420_/X 0.16fF
C4729 _385_/a_381_47# _385_/a_841_47# 0.03fF
C4730 _385_/a_558_47# _385_/a_664_47# 0.60fF
C4731 input12/a_664_47# input12/a_841_47# 0.29fF
C4732 input12/a_62_47# B[3] 0.45fF
C4733 VPWR _555_/a_382_47# 0.01fF
C4734 _455_/a_222_93# _418_/X 0.11fF
C4735 _568_/a_77_199# _568_/a_227_47# 0.24fF
C4736 _381_/C _448_/B 0.04fF
C4737 _528_/a_81_21# _527_/A 0.18fF
C4738 _528_/a_299_297# _527_/Y 0.46fF
C4739 _447_/X _628_/Y 0.77fF
C4740 _506_/Y _542_/A 0.05fF
C4741 _423_/a_215_47# _392_/Y 0.01fF
C4742 _537_/a_77_199# _537_/a_227_47# 0.24fF
C4743 _398_/a_76_199# _398_/X 0.53fF
C4744 input7/a_27_47# _489_/a_226_47# 0.00fF
C4745 _479_/a_68_297# _479_/B 0.30fF
C4746 _534_/a_209_297# _542_/B 0.00fF
C4747 _397_/X _398_/a_226_47# 0.61fF
C4748 _481_/A _376_/a_68_297# 0.30fF
C4749 _406_/A _406_/Y 0.46fF
C4750 M[13] _626_/Y 0.01fF
C4751 _471_/Y _472_/B 0.44fF
C4752 _381_/C _530_/X 0.05fF
C4753 _586_/a_76_199# _588_/A 0.02fF
C4754 _539_/A _483_/X 1.10fF
C4755 _504_/a_323_297# _627_/A 0.09fF
C4756 _557_/B _556_/A 0.02fF
C4757 _367_/a_205_297# _367_/C 0.07fF
C4758 _412_/a_226_47# _412_/a_489_413# 0.02fF
C4759 _412_/a_76_199# _412_/a_226_297# 0.01fF
C4760 _408_/B _391_/B 0.17fF
C4761 _611_/a_109_47# _610_/A 0.01fF
C4762 _563_/B _628_/Y 1.83fF
C4763 _480_/Y A[6] 0.35fF
C4764 _387_/a_78_199# _313_/A 0.43fF
C4765 _489_/X _483_/X 0.03fF
C4766 _563_/D _408_/a_68_297# 0.33fF
C4767 _433_/Y _439_/a_556_47# 0.02fF
C4768 _501_/Y _531_/C 0.31fF
C4769 _576_/a_76_199# _576_/X 0.22fF
C4770 _386_/X _518_/a_93_21# 0.21fF
C4771 _519_/A _420_/X 0.78fF
C4772 _478_/A _316_/a_381_47# 0.02fF
C4773 _447_/X _452_/X 0.18fF
C4774 B[0] _479_/a_68_297# 0.08fF
C4775 _386_/A _410_/C 0.39fF
C4776 _458_/X _458_/a_78_199# 0.21fF
C4777 _487_/a_215_47# VPWR 0.07fF
C4778 _534_/a_80_21# _535_/A 0.20fF
C4779 B[0] _541_/a_78_199# 0.17fF
C4780 _540_/a_584_47# _486_/X 0.01fF
C4781 _563_/A VPWR 6.38fF
C4782 _594_/X _574_/X 0.05fF
C4783 _520_/X _442_/D 0.03fF
C4784 _595_/X _575_/X 0.00fF
C4785 _381_/a_197_47# _381_/B 0.10fF
C4786 _513_/A _478_/a_27_47# 0.26fF
C4787 _455_/X _542_/D 0.02fF
C4788 _530_/X _570_/A 1.20fF
C4789 _520_/X _522_/a_76_199# 0.33fF
C4790 output25/a_27_47# VPWR 0.70fF
C4791 VPWR _470_/a_80_21# 0.31fF
C4792 output28/a_27_47# M[5] 0.33fF
C4793 _391_/A _392_/A 0.04fF
C4794 _516_/A A[6] 0.28fF
C4795 _542_/C _530_/X 0.05fF
C4796 A[6] _539_/A 0.18fF
C4797 _543_/B _543_/A 0.94fF
C4798 _627_/A VPWR 7.31fF
C4799 _587_/A _547_/X 0.03fF
C4800 _568_/a_227_47# _566_/A 0.15fF
C4801 _452_/A _418_/a_68_297# 0.01fF
C4802 VPWR _438_/a_68_297# 0.31fF
C4803 _556_/Y _556_/A 1.96fF
C4804 _563_/B _452_/X 0.08fF
C4805 _362_/a_489_413# _371_/B 0.13fF
C4806 _522_/a_76_199# _522_/a_489_413# 0.12fF
C4807 _404_/a_62_47# VPWR 0.71fF
C4808 _519_/X _485_/a_197_47# 0.03fF
C4809 _611_/X _591_/A 0.49fF
C4810 _533_/X _631_/Y 0.33fF
C4811 _590_/A _588_/Y 0.06fF
C4812 _455_/X _456_/X 0.60fF
C4813 _483_/a_93_21# _410_/C 0.25fF
C4814 _422_/X _421_/X 0.01fF
C4815 _554_/X _530_/X 0.03fF
C4816 _404_/a_381_47# _544_/a_558_47# 0.01fF
C4817 _543_/B _565_/a_209_47# 0.01fF
C4818 _543_/Y _565_/a_80_21# 0.31fF
C4819 _431_/X _432_/X 1.69fF
C4820 _634_/Y _374_/a_78_199# 0.01fF
C4821 _628_/a_300_47# _628_/Y 0.09fF
C4822 _338_/a_222_93# _337_/A 0.31fF
C4823 input8/a_27_47# _542_/D 0.43fF
C4824 _515_/Y _545_/Y 0.00fF
C4825 _543_/Y _545_/Y 2.61fF
C4826 VPWR _548_/X 0.89fF
C4827 _563_/a_27_297# _627_/C 0.55fF
C4828 _413_/a_68_297# _447_/B 0.47fF
C4829 _569_/A _572_/A 0.03fF
C4830 _530_/X _535_/A 1.57fF
C4831 _446_/X _457_/X 0.03fF
C4832 _492_/a_76_199# _492_/a_489_413# 0.12fF
C4833 _362_/a_226_47# VPWR 0.08fF
C4834 _469_/A _540_/X 0.03fF
C4835 _607_/a_78_199# _618_/A 0.17fF
C4836 input11/a_27_47# input3/a_62_47# 0.04fF
C4837 _573_/Y _546_/X 0.66fF
C4838 _455_/X _346_/A 1.31fF
C4839 _448_/B _419_/X 0.11fF
C4840 _340_/A _485_/D 0.15fF
C4841 _386_/A _445_/X 0.03fF
C4842 _600_/a_285_47# _601_/A 0.02fF
C4843 _567_/Y _538_/A 0.12fF
C4844 _596_/a_226_297# _616_/B 0.02fF
C4845 _413_/X _448_/B 0.43fF
C4846 _455_/X _478_/A 0.18fF
C4847 _381_/C _453_/a_93_21# 0.21fF
C4848 _565_/a_80_21# _565_/a_303_47# 0.04fF
C4849 _351_/a_27_53# VPWR 0.17fF
C4850 input5/a_558_47# input5/a_841_47# 0.07fF
C4851 _627_/D _616_/A 0.14fF
C4852 B[0] _538_/A 0.15fF
C4853 _577_/a_489_413# _576_/X 0.14fF
C4854 _577_/a_226_297# _559_/X 0.02fF
C4855 _478_/A _509_/A 0.93fF
C4856 _442_/a_109_47# VPWR 0.00fF
C4857 VPWR _368_/A 1.48fF
C4858 _327_/a_78_199# _481_/A 0.13fF
C4859 _588_/A _485_/D 0.05fF
C4860 _577_/a_76_199# _578_/a_78_199# 0.02fF
C4861 _452_/A _542_/D 1.19fF
C4862 _497_/B _496_/a_78_199# 0.21fF
C4863 output21/a_27_47# M[13] 0.43fF
C4864 _469_/a_558_47# _469_/a_664_47# 0.60fF
C4865 _598_/B _598_/A 0.93fF
C4866 VPWR _324_/a_558_47# 0.24fF
C4867 _386_/X _410_/C 0.48fF
C4868 _436_/A _421_/X 0.01fF
C4869 _566_/A _485_/D 0.18fF
C4870 _370_/a_68_297# _635_/a_300_297# 0.01fF
C4871 _330_/A _392_/A 0.37fF
C4872 _626_/Y _610_/A 0.05fF
C4873 _627_/D _572_/A 0.78fF
C4874 _468_/X _468_/a_215_47# 0.01fF
C4875 _374_/a_292_297# VPWR 0.01fF
C4876 _627_/D _622_/a_29_53# 0.65fF
C4877 _442_/A _381_/B 1.10fF
C4878 _616_/Y _624_/a_489_47# 0.16fF
C4879 output25/a_27_47# _342_/X 0.01fF
C4880 _522_/a_226_47# _521_/X 0.53fF
C4881 _588_/A _483_/X 0.00fF
C4882 _520_/X input7/a_27_47# 0.10fF
C4883 VPWR _537_/a_227_47# 0.06fF
C4884 _446_/X _503_/A 0.60fF
C4885 _608_/a_78_199# _627_/D 0.36fF
C4886 _627_/C _628_/Y 0.15fF
C4887 _445_/A _481_/A 1.01fF
C4888 _567_/B _486_/X 0.03fF
C4889 _567_/Y _488_/X 0.00fF
C4890 _442_/D _483_/a_250_297# 0.06fF
C4891 _509_/Y _631_/Y 0.35fF
C4892 _474_/Y _472_/B 0.15fF
C4893 _545_/Y _585_/B 0.21fF
C4894 _445_/A _633_/Y 0.59fF
C4895 _579_/X _602_/A 0.01fF
C4896 B[2] _612_/Y 0.03fF
C4897 _386_/a_381_47# _515_/Y 0.08fF
C4898 _444_/Y _411_/X 0.00fF
C4899 _343_/a_226_47# _343_/a_489_413# 0.02fF
C4900 _343_/a_76_199# _343_/a_226_297# 0.01fF
C4901 B[2] _390_/D 0.95fF
C4902 _627_/D _542_/D 0.55fF
C4903 _419_/a_489_413# VPWR 0.39fF
C4904 _340_/A A[6] 0.05fF
C4905 _410_/a_27_47# _442_/A 0.00fF
C4906 _455_/a_79_199# VPWR 0.67fF
C4907 _521_/a_292_297# _488_/X 0.01fF
C4908 _521_/a_493_297# _483_/X 0.02fF
C4909 M[3] A[0] 0.12fF
C4910 _505_/a_209_297# VPWR 0.45fF
C4911 _400_/a_80_21# _400_/a_209_47# 0.04fF
C4912 _583_/a_76_199# _583_/a_226_297# 0.01fF
C4913 _583_/a_226_47# _583_/a_489_413# 0.02fF
C4914 VPWR _316_/a_841_47# 0.35fF
C4915 _386_/X _445_/X 0.07fF
C4916 _498_/Y _467_/Y 0.81fF
C4917 _633_/Y _622_/C 0.03fF
C4918 VPWR _508_/a_227_47# 0.11fF
C4919 _495_/a_489_413# VPWR 0.40fF
C4920 _600_/a_27_297# B[7] 0.03fF
C4921 _577_/a_489_413# _549_/X 0.13fF
C4922 _371_/B _432_/B 0.23fF
C4923 _410_/B _410_/C 1.01fF
C4924 _378_/a_381_47# _378_/a_558_47# 0.32fF
C4925 _594_/a_27_297# _574_/a_81_21# 0.00fF
C4926 _488_/a_489_413# _559_/a_77_199# 0.05fF
C4927 _567_/B _454_/X 0.66fF
C4928 _570_/A _514_/B 0.06fF
C4929 _576_/a_226_47# _530_/X 0.06fF
C4930 _383_/X _332_/a_150_297# 0.02fF
C4931 _451_/A _541_/a_215_47# 0.06fF
C4932 _523_/X VPWR 2.08fF
C4933 _379_/a_78_199# _542_/D 0.05fF
C4934 _554_/X _556_/Y 0.01fF
C4935 _603_/Y VPWR 1.33fF
C4936 _504_/a_227_47# _468_/X 0.01fF
C4937 _542_/C _514_/B 0.39fF
C4938 _544_/A _517_/X 0.05fF
C4939 _475_/X _503_/a_558_47# 0.02fF
C4940 _419_/X _314_/a_68_297# 0.01fF
C4941 _349_/a_78_199# VPWR 0.59fF
C4942 _442_/D _503_/A 0.06fF
C4943 _417_/A _328_/A 0.21fF
C4944 _487_/a_78_199# _542_/A 0.13fF
C4945 _380_/A _381_/B 0.03fF
C4946 _614_/a_76_199# _614_/a_489_413# 0.12fF
C4947 _484_/a_215_47# _486_/A 0.01fF
C4948 _352_/a_448_47# _352_/X 0.01fF
C4949 _543_/A _451_/A 0.17fF
C4950 _396_/a_93_21# VPWR 0.37fF
C4951 _542_/A _367_/C 0.24fF
C4952 _463_/a_226_47# _463_/a_489_413# 0.02fF
C4953 _463_/a_76_199# _463_/a_226_297# 0.01fF
C4954 input12/a_62_47# _620_/a_489_413# 0.04fF
C4955 input12/a_381_47# _620_/a_226_47# 0.01fF
C4956 input12/a_558_47# _620_/a_76_199# 0.01fF
C4957 _485_/a_27_47# _547_/a_79_199# 0.04fF
C4958 _353_/X _420_/a_79_199# 0.16fF
C4959 _446_/X _471_/Y 0.96fF
C4960 _497_/B _497_/a_68_297# 0.30fF
C4961 _380_/A output28/a_27_47# 0.07fF
C4962 _360_/X _510_/A 0.03fF
C4963 _569_/Y _589_/a_489_413# 0.03fF
C4964 _469_/a_62_47# _610_/A 0.13fF
C4965 _530_/X _547_/a_544_297# 0.02fF
C4966 _442_/A _542_/A 0.63fF
C4967 _613_/a_227_297# _433_/Y 0.03fF
C4968 _579_/X _606_/A 0.06fF
C4969 _333_/a_27_47# VPWR 0.60fF
C4970 _559_/X _485_/D 0.61fF
C4971 _542_/B _385_/a_558_47# 0.02fF
C4972 _514_/B _535_/A 0.00fF
C4973 input4/a_27_47# _442_/A 0.22fF
C4974 _406_/B _631_/B 0.24fF
C4975 _613_/a_77_199# _627_/A 0.16fF
C4976 _613_/a_323_297# _612_/Y 0.01fF
C4977 _392_/Y _330_/A 0.46fF
C4978 _370_/A VPWR 1.51fF
C4979 _410_/B _445_/X 0.22fF
C4980 input3/a_381_47# _390_/D 0.61fF
C4981 _390_/D _469_/X 0.05fF
C4982 _436_/A _350_/a_27_297# 0.01fF
C4983 _386_/X _386_/A 0.96fF
C4984 _599_/Y _601_/A 0.30fF
C4985 _410_/B _584_/A 0.03fF
C4986 input5/a_62_47# _390_/B 0.14fF
C4987 _494_/a_226_47# _492_/X 0.31fF
C4988 _447_/X _447_/B 0.42fF
C4989 _557_/Y _558_/a_227_47# 0.08fF
C4990 _446_/X _446_/a_93_21# 0.13fF
C4991 M[2] _343_/a_489_413# 0.02fF
C4992 _386_/a_381_47# _386_/a_841_47# 0.03fF
C4993 _386_/a_558_47# _386_/a_664_47# 0.60fF
C4994 _447_/a_68_297# _417_/D 0.00fF
C4995 _594_/a_27_297# VPWR 0.66fF
C4996 _584_/a_68_297# _622_/X 0.20fF
C4997 _513_/A _355_/a_161_47# 0.18fF
C4998 _583_/X input12/a_664_47# 0.17fF
C4999 _446_/X _504_/X 0.22fF
C5000 _368_/B _631_/A 0.02fF
C5001 _573_/A _594_/X 0.14fF
C5002 M[7] _558_/a_323_297# 0.04fF
C5003 A[7] VPWR 1.16fF
C5004 _530_/a_226_297# _531_/B 0.02fF
C5005 _608_/a_215_47# _584_/A 0.11fF
C5006 _375_/a_544_297# _417_/A 0.04fF
C5007 _524_/a_215_47# _525_/a_226_47# 0.04fF
C5008 _367_/C _366_/a_226_47# 0.02fF
C5009 _630_/X M[5] 0.30fF
C5010 _563_/B _447_/B 0.03fF
C5011 _338_/a_222_93# VPWR 0.07fF
C5012 _386_/X _483_/a_93_21# 0.46fF
C5013 _420_/X _337_/A 0.13fF
C5014 _519_/A output32/a_27_47# 0.11fF
C5015 _614_/a_489_413# _611_/X 0.18fF
C5016 _614_/a_226_47# _613_/X 0.66fF
C5017 _550_/a_215_47# _521_/X 0.12fF
C5018 _563_/D _394_/a_62_47# 0.61fF
C5019 _575_/a_78_199# _575_/a_215_47# 0.26fF
C5020 VPWR _621_/a_215_47# 0.04fF
C5021 _600_/a_27_297# VPWR 0.89fF
C5022 _360_/X _631_/A 0.69fF
C5023 input12/a_381_47# _619_/Y 0.00fF
C5024 _376_/X _420_/a_79_199# 0.01fF
C5025 VPWR _397_/a_226_297# 0.00fF
C5026 _590_/A _592_/a_199_47# 0.07fF
C5027 _433_/Y M[6] 0.52fF
C5028 _544_/A _442_/D 0.03fF
C5029 _350_/a_27_297# _350_/X 0.20fF
C5030 _533_/a_323_297# VPWR 0.02fF
C5031 _412_/a_76_199# _419_/X 0.30fF
C5032 _587_/A _633_/Y 0.11fF
C5033 _633_/Y _612_/A 0.05fF
C5034 _326_/a_27_47# _481_/A 0.10fF
C5035 _561_/A _541_/a_215_47# 0.11fF
C5036 _380_/A _542_/A 0.32fF
C5037 _532_/a_489_47# _530_/X 0.08fF
C5038 _503_/a_664_47# VPWR 0.37fF
C5039 _410_/B _386_/A 0.47fF
C5040 _417_/D A[3] 0.05fF
C5041 _627_/A _438_/a_68_297# 0.07fF
C5042 output20/a_27_47# VPWR 0.65fF
C5043 _584_/A _395_/X 0.16fF
C5044 _493_/X _492_/X 1.82fF
C5045 _516_/a_27_47# VPWR 0.56fF
C5046 _337_/a_68_297# _631_/B 0.12fF
C5047 _334_/a_27_47# _334_/a_109_47# 0.03fF
C5048 _569_/A _570_/B 0.30fF
C5049 _569_/Y _469_/A 0.46fF
C5050 _382_/A _448_/B 0.11fF
C5051 _360_/a_76_199# _353_/X 0.31fF
C5052 _527_/B _530_/X 0.91fF
C5053 _433_/Y _547_/X 0.02fF
C5054 _597_/a_78_199# _616_/A 0.05fF
C5055 _499_/a_299_297# _497_/B 0.07fF
C5056 _390_/D _546_/X 0.04fF
C5057 _625_/Y _633_/Y 0.03fF
C5058 _436_/A _475_/A 0.39fF
C5059 _506_/Y _539_/A 0.17fF
C5060 _478_/a_27_47# VPWR 0.78fF
C5061 _313_/A _419_/X 0.01fF
C5062 _534_/a_80_21# _485_/D 0.10fF
C5063 _485_/A _520_/a_489_413# 0.02fF
C5064 _383_/a_76_199# _452_/A 0.05fF
C5065 _492_/a_76_199# _504_/X 0.02fF
C5066 _467_/Y _466_/X 0.29fF
C5067 _517_/a_68_297# _570_/A 0.33fF
C5068 _538_/Y _537_/a_227_297# 0.04fF
C5069 _490_/a_493_297# VPWR 0.01fF
C5070 _583_/X _583_/a_226_47# 0.05fF
C5071 _457_/a_489_413# VPWR 0.39fF
C5072 _540_/X _547_/X 0.04fF
C5073 _518_/a_93_21# _515_/A 0.02fF
C5074 _630_/a_76_199# _630_/a_226_47# 0.49fF
C5075 _627_/C _545_/Y 0.07fF
C5076 _544_/A _513_/a_27_47# 0.02fF
C5077 _559_/X _598_/B 0.09fF
C5078 _632_/a_215_47# _631_/B 0.16fF
C5079 _617_/a_113_297# _616_/A 0.13fF
C5080 _576_/X _574_/X 0.18fF
C5081 _335_/a_841_47# VPWR 0.32fF
C5082 _474_/Y _446_/X 0.24fF
C5083 _506_/A _410_/C 1.18fF
C5084 _490_/X _633_/Y 0.39fF
C5085 _443_/a_68_297# _346_/A 0.01fF
C5086 _570_/X _588_/A 0.57fF
C5087 _362_/a_76_199# _362_/a_489_413# 0.12fF
C5088 _509_/Y _511_/a_250_297# 0.19fF
C5089 input5/a_664_47# _431_/a_489_413# 0.03fF
C5090 input5/a_841_47# _431_/a_226_47# 0.00fF
C5091 _539_/X _472_/B 0.14fF
C5092 _566_/A _570_/X 0.17fF
C5093 _475_/a_68_297# VPWR 0.31fF
C5094 _585_/B _622_/C 0.47fF
C5095 _445_/A _359_/X 0.00fF
C5096 _476_/X _489_/X 0.19fF
C5097 _526_/a_489_413# VPWR 0.42fF
C5098 _460_/a_226_47# VPWR 0.06fF
C5099 _430_/A _371_/B 0.10fF
C5100 _328_/A _631_/B 0.20fF
C5101 _629_/A _629_/B 0.53fF
C5102 _441_/a_292_297# _340_/A 0.01fF
C5103 _426_/a_150_297# _466_/X 0.01fF
C5104 _519_/a_29_53# _519_/a_111_297# 0.01fF
C5105 _351_/A _383_/X 0.34fF
C5106 _351_/a_219_297# _351_/a_301_297# 0.02fF
C5107 _569_/A _381_/B 0.41fF
C5108 _530_/X _485_/D 1.78fF
C5109 _562_/a_78_199# _586_/S 0.03fF
C5110 _379_/a_215_47# VPWR 0.06fF
C5111 _410_/B _386_/X 0.86fF
C5112 _598_/B _616_/B 1.18fF
C5113 _493_/a_78_199# _460_/X 0.14fF
C5114 _490_/X _490_/a_215_47# 0.01fF
C5115 _625_/a_27_47# _601_/A 0.03fF
C5116 _625_/a_27_297# _624_/X 0.17fF
C5117 _527_/B _557_/B 0.12fF
C5118 _587_/A _510_/a_68_297# 0.35fF
C5119 _383_/X _397_/a_489_413# 0.00fF
C5120 _627_/C _585_/a_109_297# 0.01fF
C5121 _518_/a_346_47# _381_/B 0.04fF
C5122 _549_/a_226_47# _559_/X 0.05fF
C5123 output18/a_27_47# _558_/X 0.47fF
C5124 _406_/A _458_/a_493_297# 0.02fF
C5125 _616_/A _601_/A 0.03fF
C5126 M[2] _442_/B 0.62fF
C5127 _616_/Y _624_/X 0.90fF
C5128 _615_/a_292_297# VPWR 0.02fF
C5129 _618_/A _606_/A 2.52fF
C5130 _602_/Y _604_/a_209_297# 0.20fF
C5131 _448_/A _542_/D 0.35fF
C5132 B[1] _335_/a_664_47# 0.14fF
C5133 _349_/a_215_47# _350_/C 0.03fF
C5134 _443_/B _470_/a_209_297# 0.03fF
C5135 input12/a_841_47# VPWR 0.31fF
C5136 _466_/X _427_/A 0.82fF
C5137 _522_/X _550_/a_78_199# 0.28fF
C5138 _541_/a_215_47# VPWR 0.14fF
C5139 _327_/a_78_199# _327_/a_215_47# 0.26fF
C5140 _324_/a_381_47# _324_/a_664_47# 0.09fF
C5141 _590_/B _588_/A 0.05fF
C5142 _356_/a_292_297# _481_/A 0.02fF
C5143 _543_/Y _587_/A 0.14fF
C5144 _569_/A _469_/a_62_47# 0.13fF
C5145 _533_/X _522_/X 0.25fF
C5146 _542_/B _417_/D 0.05fF
C5147 _418_/a_68_297# _418_/A 0.30fF
C5148 _578_/a_78_199# _549_/X 0.01fF
C5149 _578_/a_215_47# _533_/X 0.18fF
C5150 _424_/a_226_297# _422_/X 0.04fF
C5151 _487_/X _472_/B 0.56fF
C5152 _563_/A _349_/a_78_199# 0.01fF
C5153 _556_/Y _527_/B 0.00fF
C5154 _623_/X _599_/Y 0.02fF
C5155 _469_/a_558_47# _586_/a_505_21# 0.00fF
C5156 _380_/A _630_/X 0.04fF
C5157 _554_/A _556_/A 0.02fF
C5158 _442_/B _332_/X 0.38fF
C5159 _502_/a_78_199# _494_/X 0.25fF
C5160 _350_/C _340_/a_27_47# 0.46fF
C5161 _633_/Y _393_/A 0.20fF
C5162 _543_/A VPWR 2.62fF
C5163 _369_/a_226_47# _343_/X 0.55fF
C5164 _544_/a_62_47# _588_/A 0.45fF
C5165 _567_/B VPWR 7.91fF
C5166 _605_/a_303_47# _602_/Y 0.02fF
C5167 _532_/a_76_199# _528_/a_81_21# 0.02fF
C5168 _386_/X _395_/X 0.43fF
C5169 _587_/A _468_/a_292_297# 0.02fF
C5170 _456_/a_76_199# _456_/a_489_413# 0.12fF
C5171 B[1] _519_/A 0.05fF
C5172 _543_/B _544_/a_841_47# 0.07fF
C5173 _631_/Y _469_/X 0.07fF
C5174 _510_/A _314_/a_68_297# 0.01fF
C5175 A[6] _530_/X 0.05fF
C5176 _444_/A _442_/D 1.15fF
C5177 _335_/a_558_47# _417_/A 0.11fF
C5178 _396_/X _400_/a_80_21# 0.00fF
C5179 _438_/X _472_/B 0.34fF
C5180 _327_/a_215_47# _445_/A 0.05fF
C5181 input9/a_27_47# _469_/A 0.10fF
C5182 _459_/a_76_199# _459_/a_226_297# 0.01fF
C5183 _363_/A VPWR 2.35fF
C5184 _500_/a_493_297# VPWR 0.01fF
C5185 _456_/X _511_/X 0.09fF
C5186 _543_/A _514_/a_150_297# 0.01fF
C5187 _520_/a_76_199# _381_/B 0.04fF
C5188 _628_/a_382_297# _628_/a_300_47# 0.02fF
C5189 _330_/A input13/a_27_47# 0.07fF
C5190 _420_/X VPWR 7.71fF
C5191 _563_/D _512_/a_215_47# 0.02fF
C5192 _429_/a_76_199# _374_/X 0.01fF
C5193 _549_/X _549_/a_76_199# 0.22fF
C5194 VPWR _468_/a_78_199# 0.59fF
C5195 _343_/a_76_199# _338_/X 0.26fF
C5196 _584_/A _394_/a_381_47# 0.61fF
C5197 _418_/A _542_/D 0.21fF
C5198 _386_/A _506_/A 0.02fF
C5199 _406_/Y _460_/X 0.40fF
C5200 _455_/a_222_93# _378_/A 0.01fF
C5201 _513_/A _485_/A 3.47fF
C5202 _511_/X _478_/A 0.03fF
C5203 _538_/A _570_/B 0.02fF
C5204 _538_/Y _469_/A 0.04fF
C5205 _382_/A _383_/a_226_47# 0.00fF
C5206 _570_/A _472_/B 0.21fF
C5207 _516_/A _359_/A 0.01fF
C5208 _436_/A _328_/B 0.08fF
C5209 _539_/a_68_297# _542_/A 0.08fF
C5210 _380_/A _363_/B 0.03fF
C5211 _587_/A _585_/B 3.19fF
C5212 _411_/A VPWR 3.65fF
C5213 B[1] _350_/a_205_297# 0.03fF
C5214 _583_/a_489_413# VPWR 0.33fF
C5215 _583_/X _581_/a_206_47# 0.05fF
C5216 _628_/a_734_297# _622_/X 0.08fF
C5217 _627_/D _593_/A 0.17fF
C5218 _519_/A _383_/X 0.03fF
C5219 _598_/B _530_/X 0.06fF
C5220 _390_/B _478_/A 0.57fF
C5221 _603_/a_27_47# _554_/X 0.06fF
C5222 _420_/X _314_/X 0.03fF
C5223 _485_/A _454_/X 0.76fF
C5224 _578_/a_292_297# _530_/X 0.08fF
C5225 _627_/a_27_297# _627_/a_205_297# 0.01fF
C5226 _411_/a_68_297# _411_/X 0.27fF
C5227 _620_/a_76_199# _618_/Y 0.34fF
C5228 _315_/a_161_47# _628_/Y 0.17fF
C5229 _430_/A _393_/A 0.22fF
C5230 _485_/A _334_/a_27_47# 0.26fF
C5231 VPWR _558_/a_77_199# 0.84fF
C5232 _410_/a_303_47# _410_/C 0.06fF
C5233 _594_/X _575_/a_215_47# 0.01fF
C5234 _506_/A _483_/a_93_21# 0.07fF
C5235 _375_/X _384_/a_76_199# 0.42fF
C5236 _613_/a_539_297# _627_/D 0.03fF
C5237 _566_/A _571_/a_346_47# 0.04fF
C5238 _456_/a_556_47# _456_/X 0.02fF
C5239 _493_/a_493_297# _457_/X 0.04fF
C5240 _505_/a_80_21# _505_/a_209_47# 0.04fF
C5241 _540_/a_256_47# _469_/X 0.06fF
C5242 _328_/X VPWR 1.32fF
C5243 _375_/a_79_199# _375_/X 0.47fF
C5244 _417_/D _563_/D 0.60fF
C5245 _591_/Y _611_/X 0.05fF
C5246 _352_/X _361_/a_226_47# 0.25fF
C5247 _570_/X _571_/a_93_21# 0.12fF
C5248 _625_/Y _585_/B 0.01fF
C5249 _469_/a_381_47# _586_/a_76_199# 0.03fF
C5250 output19/a_27_47# M[11] 0.43fF
C5251 _485_/D _514_/B 0.20fF
C5252 _448_/B _418_/B 0.77fF
C5253 _349_/a_215_47# _380_/A 0.11fF
C5254 _370_/A _368_/A 0.15fF
C5255 _408_/B _419_/X 0.86fF
C5256 _538_/Y _559_/a_227_47# 0.05fF
C5257 _583_/X _627_/B 0.18fF
C5258 _347_/A _563_/D 2.06fF
C5259 _472_/B _535_/A 0.02fF
C5260 _510_/A _385_/a_381_47# 0.12fF
C5261 _491_/X _492_/X 0.01fF
C5262 _386_/A _394_/a_381_47# 0.02fF
C5263 _469_/A _486_/X 0.99fF
C5264 _412_/a_226_47# _437_/a_79_199# 0.00fF
C5265 _412_/a_76_199# _437_/a_222_93# 0.00fF
C5266 _386_/a_664_47# VPWR 0.37fF
C5267 _627_/B _622_/X 1.55fF
C5268 input6/a_27_47# A[5] 0.41fF
C5269 _629_/A M[5] 0.12fF
C5270 _631_/B _631_/Y 0.64fF
C5271 _355_/a_161_47# VPWR 0.99fF
C5272 _422_/a_76_199# _421_/a_76_199# 0.01fF
C5273 _503_/a_664_47# _627_/A 0.05fF
C5274 VPWR _374_/X 4.91fF
C5275 _516_/A _442_/A 0.08fF
C5276 _583_/X _620_/X 1.11fF
C5277 _566_/A _546_/a_489_413# 0.11fF
C5278 _423_/a_215_47# _386_/X 0.01fF
C5279 _538_/A _381_/B 0.44fF
C5280 _386_/A _515_/A 0.69fF
C5281 _442_/A _539_/A 1.33fF
C5282 _476_/X _554_/a_68_297# 0.00fF
C5283 _342_/X _363_/A 0.01fF
C5284 _608_/X _622_/C 0.05fF
C5285 _537_/a_77_199# _537_/a_227_297# 0.13fF
C5286 _633_/Y _433_/Y 0.03fF
C5287 _386_/X _506_/A 0.19fF
C5288 _347_/A _477_/a_292_297# 0.02fF
C5289 _342_/X _420_/X 0.84fF
C5290 _351_/A _351_/a_301_297# 0.03fF
C5291 _597_/a_215_47# VPWR 0.05fF
C5292 _519_/A _484_/a_493_297# 0.02fF
C5293 _328_/X _314_/X 2.12fF
C5294 _583_/X _561_/A 0.06fF
C5295 _552_/a_226_47# _554_/A 0.05fF
C5296 _425_/a_226_47# _424_/X 0.56fF
C5297 _604_/X _557_/Y 0.18fF
C5298 _474_/A _503_/A 0.19fF
C5299 _627_/C _622_/C 2.02fF
C5300 B[0] _403_/a_27_47# 0.06fF
C5301 _554_/X _554_/A 1.60fF
C5302 _533_/a_77_199# _511_/a_250_297# 0.04fF
C5303 _334_/a_109_47# VPWR 0.01fF
C5304 VPWR _329_/X 1.81fF
C5305 _612_/A _616_/Y 0.26fF
C5306 _417_/D _518_/a_250_297# 0.14fF
C5307 _391_/A _584_/A 0.91fF
C5308 _375_/X _419_/X 0.03fF
C5309 B[7] _622_/X 0.42fF
C5310 _455_/a_448_47# _455_/X 0.01fF
C5311 _485_/A _337_/A 0.03fF
C5312 _469_/a_664_47# _584_/A 0.19fF
C5313 input13/a_27_47# _442_/B 0.29fF
C5314 _424_/X VPWR 0.14fF
C5315 _633_/Y _540_/X 0.03fF
C5316 _347_/A _518_/a_250_297# 0.06fF
C5317 _523_/a_76_199# _631_/Y 0.17fF
C5318 _385_/a_62_47# _475_/A 0.14fF
C5319 _510_/A _313_/A 0.58fF
C5320 _386_/A _385_/a_664_47# 0.05fF
C5321 _625_/Y _625_/a_27_297# 0.35fF
C5322 _553_/a_215_47# _525_/X 0.05fF
C5323 _553_/a_493_297# _524_/X 0.08fF
C5324 _569_/Y _570_/a_68_297# 0.00fF
C5325 _329_/a_489_413# _328_/X 0.14fF
C5326 VPWR _409_/a_78_199# 0.58fF
C5327 _587_/A _572_/B 0.05fF
C5328 _493_/a_78_199# _493_/X 0.21fF
C5329 input5/a_558_47# _430_/X 0.02fF
C5330 _611_/a_109_297# _622_/C 0.09fF
C5331 output31/a_27_47# _390_/B 0.26fF
C5332 _607_/X _610_/A 0.15fF
C5333 _623_/X _616_/A 0.50fF
C5334 _625_/Y _616_/Y 0.30fF
C5335 _336_/a_78_199# _442_/B 0.10fF
C5336 _426_/A _373_/Y 0.09fF
C5337 _398_/a_76_199# _399_/a_78_199# 0.04fF
C5338 _559_/X _559_/a_77_199# 0.22fF
C5339 _467_/Y _467_/a_397_297# 0.32fF
C5340 _342_/X _328_/X 0.93fF
C5341 _417_/A _447_/B 0.63fF
C5342 _627_/A _475_/a_68_297# 0.14fF
C5343 _633_/Y _610_/Y 0.12fF
C5344 _487_/X _517_/X 0.13fF
C5345 _619_/a_109_297# _619_/Y 0.05fF
C5346 _619_/a_27_47# _618_/A 0.11fF
C5347 _601_/Y _616_/Y 0.04fF
C5348 A[3] _507_/a_109_297# 0.01fF
C5349 M[8] _465_/X 0.55fF
C5350 _314_/X _329_/X 0.03fF
C5351 _475_/a_68_297# _438_/a_68_297# 0.00fF
C5352 _573_/Y _572_/A 0.14fF
C5353 M[1] VPWR 0.53fF
C5354 _612_/A _620_/a_76_199# 0.21fF
C5355 _623_/X _572_/A 0.08fF
C5356 _426_/A VPWR 2.26fF
C5357 _580_/A _390_/D 0.08fF
C5358 _327_/a_493_297# VPWR 0.02fF
C5359 _340_/A _350_/C 0.08fF
C5360 _383_/X _376_/a_150_297# 0.01fF
C5361 _602_/Y _555_/a_298_297# 0.01fF
C5362 _516_/A _380_/A 0.03fF
C5363 _623_/a_556_47# M[6] 0.02fF
C5364 _570_/X _530_/X 0.33fF
C5365 output18/a_27_47# _501_/a_397_297# 0.01fF
C5366 _473_/a_539_297# VPWR 0.02fF
C5367 _382_/B _420_/a_79_199# 0.22fF
C5368 _590_/B _592_/a_113_297# 0.09fF
C5369 _386_/X _515_/A 1.38fF
C5370 _626_/Y _511_/X 1.01fF
C5371 _480_/A _505_/a_80_21# 0.02fF
C5372 M[13] _626_/a_109_47# 0.00fF
C5373 _476_/a_250_297# _587_/A 0.02fF
C5374 _369_/a_226_47# _370_/B 0.05fF
C5375 _381_/C _517_/X 0.06fF
C5376 _584_/A A[3] 0.09fF
C5377 _416_/a_78_199# M[9] 0.03fF
C5378 _329_/a_489_413# _329_/X 0.00fF
C5379 _474_/A _471_/Y 1.19fF
C5380 _604_/X _606_/A 0.02fF
C5381 _545_/Y _469_/X 1.12fF
C5382 _563_/A _541_/a_215_47# 0.01fF
C5383 _513_/A _383_/X 0.11fF
C5384 _420_/a_222_93# _452_/A 0.00fF
C5385 _628_/a_28_47# VPWR 0.10fF
C5386 _441_/a_493_297# _346_/A 0.11fF
C5387 _370_/a_68_297# _370_/B 0.30fF
C5388 _504_/a_77_199# _478_/A 0.17fF
C5389 _626_/Y _390_/B 0.27fF
C5390 _626_/Y _601_/A 0.25fF
C5391 _347_/A _518_/X 0.03fF
C5392 _493_/X _626_/Y 0.24fF
C5393 _340_/A _442_/A 0.21fF
C5394 _476_/a_93_21# VPWR 0.17fF
C5395 _519_/X _547_/a_448_47# 0.15fF
C5396 _628_/a_300_47# _625_/Y 0.09fF
C5397 _540_/a_93_21# _472_/B 0.15fF
C5398 _342_/X _329_/X 0.11fF
C5399 _589_/a_226_47# _589_/a_489_413# 0.02fF
C5400 _589_/a_76_199# _589_/a_226_297# 0.01fF
C5401 _511_/a_250_297# _469_/X 0.06fF
C5402 _505_/a_80_21# _481_/A 0.10fF
C5403 _408_/a_68_297# _394_/a_558_47# 0.01fF
C5404 M[0] _631_/Y 0.10fF
C5405 _565_/a_80_21# _512_/a_78_199# 0.02fF
C5406 _350_/a_277_297# _563_/A 0.03fF
C5407 _419_/X _458_/a_215_47# 0.23fF
C5408 _465_/a_109_297# _465_/X 0.03fF
C5409 _612_/Y _599_/Y 0.09fF
C5410 _474_/Y _476_/a_584_47# 0.01fF
C5411 _374_/X _399_/a_215_47# 0.11fF
C5412 _581_/B _530_/X 0.10fF
C5413 _571_/a_93_21# _571_/a_346_47# 0.05fF
C5414 _517_/X _570_/A 1.26fF
C5415 _454_/X _383_/X 0.23fF
C5416 _452_/a_68_297# _628_/Y 0.22fF
C5417 VPWR _553_/a_78_199# 0.63fF
C5418 _429_/a_76_199# _429_/a_226_47# 0.49fF
C5419 _633_/Y _443_/B 0.01fF
C5420 M[8] M[10] 0.03fF
C5421 _417_/A _343_/X 0.27fF
C5422 _583_/X VPWR 4.88fF
C5423 _499_/a_81_21# _498_/Y 0.48fF
C5424 _390_/B _406_/Y 0.10fF
C5425 input3/a_664_47# _485_/D 0.12fF
C5426 _563_/D _477_/a_78_199# 0.17fF
C5427 _626_/Y _549_/a_489_413# 0.09fF
C5428 _595_/a_539_297# VPWR 0.02fF
C5429 VPWR _622_/X 2.01fF
C5430 _587_/A _509_/Y 0.15fF
C5431 _543_/A _627_/A 0.13fF
C5432 _440_/X _457_/X 0.69fF
C5433 _567_/B _627_/A 0.05fF
C5434 _384_/X _350_/X 0.12fF
C5435 _574_/a_81_21# _574_/a_299_297# 0.21fF
C5436 _422_/a_76_199# _422_/a_226_47# 0.49fF
C5437 _570_/B _595_/a_77_199# 0.01fF
C5438 _567_/Y _390_/D 0.25fF
C5439 _629_/A _630_/a_226_297# 0.02fF
C5440 _537_/a_227_297# VPWR 0.01fF
C5441 _370_/a_68_297# _371_/B 0.27fF
C5442 B[1] _337_/A 0.02fF
C5443 _567_/B _438_/a_68_297# 0.00fF
C5444 _390_/D B[0] 0.05fF
C5445 _627_/C _612_/A 0.44fF
C5446 _404_/a_62_47# _543_/A 0.07fF
C5447 _442_/B _410_/C 0.12fF
C5448 _382_/a_68_297# _382_/X 0.28fF
C5449 _500_/a_78_199# _464_/A 0.15fF
C5450 _542_/A _488_/X 0.08fF
C5451 _542_/B _410_/C 1.29fF
C5452 _487_/X _442_/D 0.03fF
C5453 VPWR _369_/a_76_199# 0.45fF
C5454 _423_/X _393_/A 0.19fF
C5455 _411_/B _475_/A 0.19fF
C5456 _543_/B _547_/X 0.01fF
C5457 _477_/a_78_199# _477_/a_292_297# 0.03fF
C5458 _563_/D _518_/a_93_21# 0.12fF
C5459 _519_/X _520_/a_76_199# 0.25fF
C5460 VPWR output32/a_27_47# 0.74fF
C5461 _417_/D _520_/X 0.08fF
C5462 _452_/a_68_297# _452_/X 0.27fF
C5463 _525_/a_76_199# _525_/a_226_47# 0.49fF
C5464 _627_/A _468_/a_78_199# 0.00fF
C5465 _511_/a_584_47# _433_/Y 0.03fF
C5466 _347_/A _520_/X 0.10fF
C5467 _625_/Y _627_/C 0.22fF
C5468 _580_/a_68_297# VPWR 0.31fF
C5469 _337_/B _419_/X 0.36fF
C5470 _516_/A _455_/X 0.92fF
C5471 _455_/X _539_/A 0.16fF
C5472 _475_/X VPWR 1.29fF
C5473 _373_/a_113_297# _629_/B 0.09fF
C5474 _411_/A _470_/a_80_21# 0.10fF
C5475 _422_/X _406_/B 0.26fF
C5476 _440_/X _459_/X 1.91fF
C5477 _589_/a_226_297# _612_/A 0.04fF
C5478 _610_/A _588_/A 0.80fF
C5479 _483_/a_346_47# _542_/A 0.02fF
C5480 _477_/a_78_199# _518_/a_250_297# 0.02fF
C5481 _429_/a_489_413# _371_/B 0.13fF
C5482 input10/a_27_47# _350_/X 0.02fF
C5483 _469_/A B[7] 0.02fF
C5484 _545_/Y _546_/X 0.18fF
C5485 _631_/a_109_297# _631_/B 0.01fF
C5486 _493_/X _527_/A 0.01fF
C5487 _539_/A _509_/A 0.18fF
C5488 B[2] _624_/X 0.01fF
C5489 _469_/a_558_47# _503_/A 0.05fF
C5490 _336_/a_78_199# _336_/a_292_297# 0.03fF
C5491 _562_/a_78_199# _564_/A 0.21fF
C5492 _426_/A _399_/a_215_47# 0.01fF
C5493 _602_/A _554_/B 0.03fF
C5494 _337_/A _383_/X 0.40fF
C5495 _391_/B _394_/a_62_47# 0.15fF
C5496 _589_/a_489_413# VPWR 0.39fF
C5497 _376_/X _383_/a_226_297# 0.03fF
C5498 _412_/X _458_/X 0.13fF
C5499 _445_/X _442_/B 0.05fF
C5500 _585_/B _433_/Y 0.21fF
C5501 _534_/a_209_47# _515_/A 0.06fF
C5502 _430_/X _466_/X 0.02fF
C5503 _626_/Y _524_/X 0.10fF
C5504 _542_/B _445_/X 0.17fF
C5505 _475_/A _366_/a_226_47# 0.00fF
C5506 _396_/X _397_/a_489_413# 0.16fF
C5507 _429_/a_226_47# VPWR 0.07fF
C5508 _487_/X _521_/a_215_47# 0.10fF
C5509 _584_/A _442_/B 1.44fF
C5510 _448_/A _542_/A 0.78fF
C5511 _556_/A _558_/a_227_47# 0.16fF
C5512 VPWR _574_/a_299_297# 0.67fF
C5513 _442_/D _570_/A 0.03fF
C5514 _538_/Y _570_/a_68_297# 0.00fF
C5515 _459_/a_226_47# _458_/X 0.52fF
C5516 _563_/B _484_/a_78_199# 0.13fF
C5517 _518_/a_93_21# _518_/a_250_297# 0.50fF
C5518 _442_/D _316_/a_62_47# 0.00fF
C5519 _504_/a_227_47# _587_/A 0.02fF
C5520 _437_/a_448_47# _411_/X 0.24fF
C5521 _596_/a_226_297# _594_/X 0.03fF
C5522 _596_/a_489_413# _595_/X 0.14fF
C5523 _485_/A VPWR 4.10fF
C5524 _542_/C _442_/D 0.81fF
C5525 _430_/A _365_/a_299_297# 0.02fF
C5526 _360_/X _350_/C 0.83fF
C5527 output25/a_27_47# _374_/X 0.00fF
C5528 _368_/B _367_/C 0.15fF
C5529 _423_/a_78_199# _384_/X 0.42fF
C5530 _408_/B _510_/A 0.91fF
C5531 _417_/A _350_/B 0.02fF
C5532 _605_/a_209_297# _557_/B 0.00fF
C5533 _474_/A _474_/Y 0.72fF
C5534 _386_/X _330_/A 1.39fF
C5535 _504_/a_539_297# VPWR 0.02fF
C5536 _634_/Y VPWR 1.67fF
C5537 _425_/a_226_47# _425_/a_489_413# 0.02fF
C5538 _425_/a_76_199# _425_/a_226_297# 0.01fF
C5539 _322_/A _347_/A 0.11fF
C5540 _596_/a_76_199# _596_/a_226_297# 0.01fF
C5541 _596_/a_226_47# _596_/a_489_413# 0.02fF
C5542 _342_/X _369_/a_76_199# 0.39fF
C5543 _516_/A _477_/a_215_47# 0.27fF
C5544 _563_/D _410_/C 0.87fF
C5545 _516_/A _452_/A 0.33fF
C5546 _613_/X A[3] 0.15fF
C5547 _503_/a_558_47# _503_/a_841_47# 0.07fF
C5548 _350_/C _409_/a_215_47# 0.07fF
C5549 _353_/X _382_/B 0.54fF
C5550 _569_/A _435_/a_27_47# 0.07fF
C5551 _547_/X _486_/X 0.12fF
C5552 _563_/A _334_/a_109_47# 0.03fF
C5553 _554_/X _579_/X 0.22fF
C5554 B[2] _618_/Y 0.02fF
C5555 _392_/A _391_/B 0.01fF
C5556 _442_/D _535_/A 0.03fF
C5557 _593_/A _601_/A 0.38fF
C5558 _367_/a_27_297# VPWR 0.30fF
C5559 _510_/A _472_/B 2.72fF
C5560 _547_/a_79_199# _547_/a_222_93# 0.51fF
C5561 _513_/A _547_/X 0.38fF
C5562 _585_/B _610_/Y 0.01fF
C5563 _425_/a_489_413# VPWR 0.33fF
C5564 _328_/A _352_/X 0.02fF
C5565 _418_/B _378_/a_62_47# 0.12fF
C5566 _360_/X _442_/A 0.02fF
C5567 _411_/B _390_/B 0.12fF
C5568 _578_/a_215_47# _551_/a_226_47# 0.02fF
C5569 VPWR _501_/a_109_297# 0.01fF
C5570 _536_/Y _538_/A 0.00fF
C5571 _563_/A _409_/a_78_199# 0.01fF
C5572 _423_/X _433_/Y 0.03fF
C5573 _467_/Y _498_/A 0.16fF
C5574 _612_/Y _625_/a_27_47# 0.24fF
C5575 output18/a_27_47# _531_/A 0.01fF
C5576 _539_/a_68_297# _539_/A 0.39fF
C5577 _487_/a_493_297# _563_/B 0.01fF
C5578 _386_/A _442_/B 2.09fF
C5579 _542_/B _386_/A 0.98fF
C5580 _574_/X _575_/a_292_297# 0.02fF
C5581 _605_/a_80_21# _604_/X 0.35fF
C5582 _605_/a_209_297# _556_/Y 0.22fF
C5583 _440_/a_76_199# _436_/X 0.17fF
C5584 _518_/a_93_21# _518_/X 0.13fF
C5585 _375_/X _510_/A 0.17fF
C5586 _455_/X _340_/A 0.03fF
C5587 _612_/Y _616_/A 0.25fF
C5588 _513_/a_109_47# _542_/B 0.01fF
C5589 _539_/A _540_/a_250_297# 0.20fF
C5590 _338_/X _337_/B 0.38fF
C5591 _436_/a_150_297# _436_/a_68_297# 0.02fF
C5592 _513_/a_27_47# _542_/C 0.23fF
C5593 _544_/a_841_47# VPWR 0.32fF
C5594 _469_/A VPWR 2.61fF
C5595 B[0] _563_/a_27_297# 0.11fF
C5596 _586_/S _563_/B 0.01fF
C5597 _408_/B _631_/A 0.12fF
C5598 _391_/A _395_/X 0.11fF
C5599 _594_/a_109_297# _615_/a_78_199# 0.01fF
C5600 _524_/a_78_199# _490_/X 0.13fF
C5601 _493_/X _502_/a_493_297# 0.08fF
C5602 _381_/C _358_/a_27_47# 0.19fF
C5603 _365_/a_384_47# _363_/A 0.09fF
C5604 _544_/a_664_47# _544_/a_841_47# 0.29fF
C5605 _563_/D _445_/X 0.74fF
C5606 _518_/X _547_/a_79_199# 0.03fF
C5607 _623_/X _626_/Y 0.38fF
C5608 _488_/a_76_199# _486_/X 0.41fF
C5609 _498_/Y _497_/A 0.52fF
C5610 _599_/A VPWR 2.19fF
C5611 _374_/a_292_297# _374_/X 0.02fF
C5612 _563_/D _584_/A 1.47fF
C5613 _483_/X _472_/B 0.06fF
C5614 _335_/a_664_47# _633_/Y 0.08fF
C5615 _431_/a_76_199# _428_/X 0.44fF
C5616 _431_/a_226_47# _430_/X 0.53fF
C5617 _544_/A _378_/a_381_47# 0.61fF
C5618 _613_/a_77_199# _622_/X 0.02fF
C5619 _624_/a_76_199# _624_/a_206_369# 0.69fF
C5620 _622_/C _469_/X 0.86fF
C5621 _376_/X _382_/B 0.05fF
C5622 _569_/A _568_/a_77_199# 0.24fF
C5623 _606_/Y _599_/A 0.10fF
C5624 _577_/a_226_47# _577_/a_489_413# 0.02fF
C5625 _577_/a_76_199# _577_/a_226_297# 0.01fF
C5626 _417_/D _503_/A 0.05fF
C5627 _390_/B _470_/a_303_47# 0.03fF
C5628 _516_/A _379_/a_78_199# 0.13fF
C5629 VPWR _559_/a_227_47# 0.05fF
C5630 _491_/X _626_/Y 0.41fF
C5631 _635_/Y M[3] 0.06fF
C5632 _564_/a_219_297# _621_/X 0.01fF
C5633 _480_/Y _479_/a_68_297# 0.01fF
C5634 _458_/X _631_/B 0.19fF
C5635 B[1] VPWR 4.56fF
C5636 _610_/A _616_/B 0.11fF
C5637 _610_/Y _616_/Y 0.16fF
C5638 _378_/A _447_/X 0.03fF
C5639 _516_/A _520_/a_76_199# 0.15fF
C5640 VPWR _489_/a_76_199# 0.53fF
C5641 _375_/a_448_47# _359_/X 0.14fF
C5642 _628_/a_300_47# _586_/S 0.00fF
C5643 _375_/X _631_/A 1.32fF
C5644 _360_/X _380_/A 0.01fF
C5645 _519_/A _481_/A 0.14fF
C5646 _436_/A _332_/a_68_297# 0.33fF
C5647 B[0] _628_/Y 0.03fF
C5648 _447_/a_68_297# M[9] 0.07fF
C5649 _477_/a_215_47# _479_/A 0.01fF
C5650 _633_/Y _519_/A 0.03fF
C5651 _542_/B _386_/X 0.03fF
C5652 A[6] _472_/B 0.05fF
C5653 _587_/A _533_/a_77_199# 0.02fF
C5654 _340_/A _477_/a_215_47# 0.07fF
C5655 _613_/a_227_297# B[7] 0.04fF
C5656 _520_/X _518_/a_93_21# 0.07fF
C5657 _476_/a_93_21# _627_/A 0.01fF
C5658 _584_/A _586_/a_505_21# 0.12fF
C5659 _525_/a_226_47# _492_/a_226_47# 0.00fF
C5660 _525_/a_489_413# _492_/a_76_199# 0.02fF
C5661 B[2] _612_/A 0.43fF
C5662 _516_/A _479_/a_68_297# 0.02fF
C5663 _330_/A _395_/X 0.34fF
C5664 _394_/a_62_47# _394_/a_558_47# 0.03fF
C5665 _479_/a_68_297# _539_/A 0.01fF
C5666 _392_/Y _391_/B 0.10fF
C5667 _496_/a_78_199# _462_/X 0.30fF
C5668 _460_/X _462_/a_226_47# 0.31fF
C5669 _381_/C _359_/B 0.04fF
C5670 _386_/A _563_/D 0.17fF
C5671 B[7] output23/a_27_47# 0.10fF
C5672 _378_/A _563_/B 0.30fF
C5673 _468_/X _492_/X 0.59fF
C5674 M[6] _627_/B 0.43fF
C5675 _562_/a_215_47# _451_/a_27_47# 0.03fF
C5676 _349_/a_215_47# _475_/A 0.05fF
C5677 _504_/X _554_/B 0.19fF
C5678 _360_/a_489_413# _375_/X 0.01fF
C5679 _448_/B _367_/C 0.66fF
C5680 _460_/a_76_199# _460_/a_489_413# 0.12fF
C5681 _569_/A _588_/A 2.04fF
C5682 _627_/A _595_/a_539_297# 0.03fF
C5683 VPWR _466_/a_493_297# 0.01fF
C5684 _408_/X _631_/Y 0.15fF
C5685 _523_/a_76_199# _522_/X 0.23fF
C5686 _523_/a_226_47# _511_/X 0.24fF
C5687 _465_/a_373_47# _465_/a_27_297# 0.08fF
C5688 _385_/a_381_47# _388_/a_27_47# 0.04fF
C5689 _383_/X VPWR 4.12fF
C5690 B[2] _625_/Y 0.09fF
C5691 _569_/A _566_/A 0.56fF
C5692 _485_/a_303_47# _542_/A 0.03fF
C5693 _390_/D _478_/A 0.03fF
C5694 _608_/X _586_/S 0.25fF
C5695 _329_/a_226_297# _314_/X 0.01fF
C5696 _356_/a_215_47# VPWR 0.06fF
C5697 _509_/Y _433_/Y 0.70fF
C5698 _442_/D _621_/X 0.76fF
C5699 _612_/Y _619_/Y 0.08fF
C5700 _454_/a_226_47# _628_/Y 0.06fF
C5701 _382_/X _320_/a_161_47# 0.00fF
C5702 _375_/a_79_199# _359_/B 0.19fF
C5703 _631_/B _350_/B 0.16fF
C5704 _627_/C _433_/Y 0.02fF
C5705 B[0] _481_/a_27_47# 0.06fF
C5706 _405_/a_109_297# VPWR 0.01fF
C5707 _425_/a_226_47# _407_/Y 0.22fF
C5708 output21/a_27_47# _623_/X 0.00fF
C5709 _355_/A _479_/B 0.14fF
C5710 _627_/C _586_/S 1.86fF
C5711 _544_/A _417_/D 0.37fF
C5712 _385_/a_381_47# _394_/a_664_47# 0.01fF
C5713 _410_/B _442_/B 0.03fF
C5714 _627_/D _588_/A 0.49fF
C5715 _410_/B _542_/B 0.44fF
C5716 _532_/a_206_369# _532_/a_489_47# 0.04fF
C5717 _428_/a_384_47# _426_/A 0.10fF
C5718 _475_/X _627_/A 0.38fF
C5719 _544_/A _347_/A 0.35fF
C5720 _475_/X _438_/a_68_297# 0.01fF
C5721 _584_/A _518_/X 0.03fF
C5722 B[0] _540_/a_256_47# 0.01fF
C5723 _510_/X _539_/A 0.18fF
C5724 _510_/A _337_/B 0.01fF
C5725 _580_/A _579_/a_145_75# 0.02fF
C5726 _459_/a_76_199# VPWR 0.51fF
C5727 _527_/B _532_/a_206_369# 0.42fF
C5728 _407_/Y VPWR 1.68fF
C5729 _599_/Y _624_/a_489_47# 0.12fF
C5730 _612_/Y _589_/a_556_47# 0.02fF
C5731 _587_/A _469_/X 1.76fF
C5732 _360_/X _455_/X 0.36fF
C5733 _519_/C _453_/a_250_297# 0.12fF
C5734 _370_/A _329_/X 0.01fF
C5735 VPWR _484_/a_493_297# 0.01fF
C5736 _519_/A _413_/a_68_297# 0.03fF
C5737 _386_/X _563_/D 0.56fF
C5738 _563_/A _485_/A 0.72fF
C5739 _480_/A _486_/X 0.78fF
C5740 _346_/a_161_47# _322_/a_27_47# 0.03fF
C5741 _573_/Y _593_/A 0.69fF
C5742 _573_/A _593_/Y 0.46fF
C5743 _419_/X _408_/a_68_297# 0.01fF
C5744 _329_/a_226_47# _417_/A 0.06fF
C5745 _569_/Y _585_/B 0.03fF
C5746 _386_/a_558_47# _480_/A 0.02fF
C5747 _386_/a_62_47# _480_/Y 0.02fF
C5748 _613_/a_227_297# VPWR 0.01fF
C5749 _627_/C _610_/Y 0.16fF
C5750 _385_/a_558_47# _385_/a_841_47# 0.07fF
C5751 _562_/a_78_199# _627_/B 0.25fF
C5752 input12/a_62_47# _442_/D 0.31fF
C5753 input12/a_381_47# B[3] 0.02fF
C5754 input3/a_62_47# VPWR 0.53fF
C5755 _517_/X _485_/D 0.02fF
C5756 _510_/A _446_/X 0.03fF
C5757 _455_/a_544_297# _418_/X 0.06fF
C5758 _551_/a_76_199# VPWR 0.49fF
C5759 _611_/a_27_297# _633_/Y 0.14fF
C5760 _453_/X _628_/Y 0.15fF
C5761 _423_/a_215_47# _330_/A 0.01fF
C5762 _528_/a_299_297# _527_/A 0.12fF
C5763 _623_/X _613_/a_539_297# 0.02fF
C5764 _398_/a_226_47# _398_/X 0.20fF
C5765 _497_/a_68_297# _462_/X 0.01fF
C5766 _479_/a_68_297# _479_/A 0.32fF
C5767 output25/a_27_47# _634_/Y 0.48fF
C5768 _406_/B _406_/Y 0.47fF
C5769 _541_/a_78_199# _340_/A 0.42fF
C5770 _397_/X _398_/a_489_413# 0.14fF
C5771 _547_/X _574_/a_81_21# 0.06fF
C5772 _472_/Y _472_/B 1.09fF
C5773 _318_/a_27_47# _410_/C 0.29fF
C5774 VPWR output23/a_27_47# 0.80fF
C5775 _466_/a_78_199# _466_/a_215_47# 0.26fF
C5776 input11/a_27_47# B[2] 0.38fF
C5777 _481_/A _486_/X 0.68fF
C5778 _436_/X _438_/X 0.04fF
C5779 _504_/a_539_297# _627_/A 0.03fF
C5780 _502_/a_78_199# VPWR 0.77fF
C5781 _338_/X _344_/a_493_297# 0.08fF
C5782 _380_/A _530_/X 0.05fF
C5783 _563_/a_27_297# _542_/D 0.25fF
C5784 _532_/a_489_47# _498_/Y 0.12fF
C5785 _378_/A _627_/C 0.14fF
C5786 _516_/A _386_/a_62_47# 0.14fF
C5787 _633_/Y _486_/X 0.01fF
C5788 _367_/a_277_297# _367_/C 0.01fF
C5789 _513_/A _481_/A 0.62fF
C5790 _611_/a_373_47# _610_/A 0.01fF
C5791 _387_/a_292_297# _313_/A 0.01fF
C5792 _489_/X _488_/X 0.01fF
C5793 _543_/A _541_/a_215_47# 0.01fF
C5794 _527_/B _498_/Y 0.02fF
C5795 _444_/Y _411_/B 0.19fF
C5796 _520_/X _584_/A 0.08fF
C5797 _491_/a_489_413# _633_/Y 0.09fF
C5798 _576_/a_76_199# _575_/X 0.22fF
C5799 _576_/a_226_47# _576_/X 0.05fF
C5800 _386_/X _518_/a_250_297# 0.03fF
C5801 _360_/X B[4] 0.01fF
C5802 _453_/X _452_/X 0.40fF
C5803 _523_/X _553_/a_78_199# 0.01fF
C5804 _603_/Y _553_/a_78_199# 0.11fF
C5805 _534_/a_209_297# _535_/A 0.04fF
C5806 _584_/A _590_/A 0.07fF
C5807 _491_/a_76_199# _489_/X 0.47fF
C5808 _342_/a_68_297# _350_/C 0.30fF
C5809 _410_/B _563_/D 0.03fF
C5810 _390_/B _340_/a_27_47# 0.10fF
C5811 _420_/a_79_199# _420_/a_448_47# 0.13fF
C5812 _440_/a_76_199# _440_/X 0.22fF
C5813 _520_/X _522_/a_226_47# 0.28fF
C5814 _454_/X _481_/A 0.83fF
C5815 VPWR _470_/a_209_297# 0.45fF
C5816 VPWR M[6] 1.27fF
C5817 _349_/a_493_297# _350_/B 0.04fF
C5818 _543_/B _543_/Y 1.35fF
C5819 _633_/Y _454_/X 0.23fF
C5820 _604_/X _556_/A 0.34fF
C5821 _587_/A _546_/X 0.03fF
C5822 _596_/a_76_199# _598_/B 0.02fF
C5823 _330_/A _361_/X 0.39fF
C5824 _634_/Y _368_/A 0.75fF
C5825 _469_/A _627_/A 0.83fF
C5826 A[6] _517_/X 0.32fF
C5827 _626_/Y _612_/Y 0.03fF
C5828 _530_/X _552_/a_489_413# 0.09fF
C5829 _522_/a_76_199# _522_/a_226_297# 0.01fF
C5830 _522_/a_226_47# _522_/a_489_413# 0.02fF
C5831 _404_/a_381_47# VPWR 0.42fF
C5832 _390_/D _626_/Y 0.03fF
C5833 _436_/A _631_/Y 0.03fF
C5834 _483_/a_250_297# _410_/C 0.18fF
C5835 _611_/X _621_/X 0.01fF
C5836 _613_/X _591_/A 1.03fF
C5837 _542_/D _628_/Y 0.09fF
C5838 _543_/B _565_/a_303_47# 0.01fF
C5839 _543_/Y _565_/a_209_297# 0.09fF
C5840 _531_/B _531_/a_109_297# 0.07fF
C5841 _404_/a_381_47# _544_/a_664_47# 0.04fF
C5842 _431_/X _430_/X 0.22fF
C5843 _569_/A _571_/a_93_21# 0.46fF
C5844 _338_/a_544_297# _337_/A 0.01fF
C5845 VPWR _547_/X 14.19fF
C5846 _442_/D _485_/D 0.03fF
C5847 _417_/a_197_47# _542_/A 0.03fF
C5848 _413_/a_150_297# _447_/B 0.02fF
C5849 _490_/a_215_47# _454_/X 0.41fF
C5850 _563_/a_109_297# _627_/C 0.04fF
C5851 _362_/a_489_413# VPWR 0.39fF
C5852 _357_/a_27_47# _478_/A 0.40fF
C5853 _567_/B _468_/a_78_199# 0.18fF
C5854 _492_/a_76_199# _492_/a_226_297# 0.01fF
C5855 _492_/a_226_47# _492_/a_489_413# 0.02fF
C5856 _603_/a_27_47# _581_/B 0.03fF
C5857 _437_/X _472_/B 0.15fF
C5858 A[1] VPWR 0.38fF
C5859 M[2] B[5] 0.05fF
C5860 _368_/a_68_297# VPWR 0.29fF
C5861 _455_/X _448_/B 1.08fF
C5862 B[1] _563_/A 1.38fF
C5863 _386_/A _520_/X 0.86fF
C5864 _381_/C _453_/a_250_297# 0.06fF
C5865 VPWR _570_/a_68_297# 0.30fF
C5866 _322_/A _584_/A 0.85fF
C5867 input5/a_62_47# A[4] 0.45fF
C5868 input5/a_664_47# input5/a_841_47# 0.29fF
C5869 _386_/X _518_/X 0.03fF
C5870 _359_/X _519_/A 0.03fF
C5871 _468_/X _478_/A 0.09fF
C5872 A[3] _535_/Y 0.03fF
C5873 _511_/X _539_/A 0.40fF
C5874 _442_/a_197_47# VPWR 0.00fF
C5875 _382_/X _542_/D 0.26fF
C5876 _544_/A _477_/a_78_199# 0.33fF
C5877 M[11] _628_/Y 0.00fF
C5878 _452_/X _542_/D 0.64fF
C5879 _437_/a_448_47# _408_/X 0.14fF
C5880 output27/a_27_47# _373_/Y 0.45fF
C5881 _348_/a_27_47# VPWR 0.69fF
C5882 VPWR _324_/a_664_47# 0.37fF
C5883 _520_/X _521_/X 1.80fF
C5884 _456_/X _631_/Y 0.12fF
C5885 _381_/B _486_/A 0.13fF
C5886 _629_/X VPWR 0.95fF
C5887 _429_/a_76_199# _432_/B 0.22fF
C5888 _511_/X _489_/X 0.05fF
C5889 _607_/X _601_/A 1.08fF
C5890 _542_/B _506_/A 0.38fF
C5891 _585_/B _507_/Y 0.63fF
C5892 _374_/a_493_297# VPWR 0.01fF
C5893 _543_/B _585_/B 0.25fF
C5894 _313_/A _350_/C 0.47fF
C5895 _627_/D _622_/a_111_297# 0.01fF
C5896 _463_/a_76_199# _497_/a_68_297# 0.00fF
C5897 _381_/a_27_47# _382_/B 0.18fF
C5898 _330_/A input1/a_27_47# 0.22fF
C5899 _616_/B _624_/a_205_47# 0.08fF
C5900 output27/a_27_47# VPWR 0.70fF
C5901 _598_/A _601_/A 0.32fF
C5902 _390_/D _381_/B 0.05fF
C5903 _439_/a_76_199# _436_/a_68_297# 0.01fF
C5904 _488_/a_76_199# VPWR 0.51fF
C5905 _447_/X _519_/A 1.24fF
C5906 _522_/a_489_413# _521_/X 0.17fF
C5907 _562_/a_78_199# VPWR 0.64fF
C5908 _529_/a_27_47# _531_/A 0.11fF
C5909 _631_/Y _478_/A 0.18fF
C5910 _484_/a_78_199# _484_/a_215_47# 0.26fF
C5911 _352_/a_79_199# _352_/a_222_93# 0.51fF
C5912 _608_/a_292_297# _627_/D 0.08fF
C5913 _515_/Y _486_/X 0.06fF
C5914 _557_/A _557_/a_109_297# 0.01fF
C5915 _449_/A _519_/C 1.66fF
C5916 _442_/D _483_/a_256_47# 0.03fF
C5917 _544_/A _547_/a_79_199# 0.07fF
C5918 _458_/X _460_/a_226_297# 0.02fF
C5919 _328_/B _328_/a_68_297# 0.30fF
C5920 _506_/Y _472_/B 0.26fF
C5921 A[6] _442_/D 0.05fF
C5922 _386_/a_558_47# _515_/Y 0.10fF
C5923 _513_/A _543_/Y 1.35fF
C5924 _420_/X _328_/X 0.53fF
C5925 _591_/A _590_/a_68_297# 0.27fF
C5926 _569_/Y _595_/a_227_47# 0.07fF
C5927 _448_/B _452_/A 0.29fF
C5928 _586_/a_218_374# _588_/A 0.02fF
C5929 _455_/a_222_93# VPWR 0.07fF
C5930 _400_/a_80_21# _400_/a_303_47# 0.04fF
C5931 _563_/B _519_/A 0.55fF
C5932 _521_/a_493_297# _488_/X 0.03fF
C5933 _521_/a_78_199# _486_/X 0.01fF
C5934 _521_/a_215_47# _483_/X 0.15fF
C5935 _613_/a_77_199# _613_/a_227_297# 0.13fF
C5936 _566_/Y _595_/X 0.15fF
C5937 _386_/X _520_/X 0.91fF
C5938 _495_/a_226_297# VPWR 0.00fF
C5939 _442_/B _361_/X 0.17fF
C5940 _600_/a_114_47# B[7] 0.05fF
C5941 _359_/a_68_297# _359_/a_150_297# 0.02fF
C5942 _580_/A _578_/a_215_47# 0.08fF
C5943 _378_/a_381_47# _378_/a_664_47# 0.09fF
C5944 _476_/X _472_/B 0.28fF
C5945 _390_/a_27_47# _410_/C 0.15fF
C5946 _386_/X _437_/a_79_199# 0.02fF
C5947 _442_/B _394_/a_381_47# 0.12fF
C5948 _347_/A _387_/a_78_199# 0.01fF
C5949 _576_/a_489_413# _530_/X 0.11fF
C5950 _569_/Y _627_/C 0.03fF
C5951 _456_/X _490_/a_78_199# 0.36fF
C5952 _520_/X _550_/a_215_47# 0.16fF
C5953 _457_/a_76_199# _456_/X 0.21fF
C5954 _634_/Y _370_/A 0.54fF
C5955 VPWR _432_/B 1.62fF
C5956 _584_/A _503_/A 0.70fF
C5957 _432_/A _629_/A 0.38fF
C5958 _542_/B _515_/A 0.65fF
C5959 _619_/Y _607_/a_215_47# 0.02fF
C5960 _475_/X _503_/a_664_47# 0.02fF
C5961 _417_/A _351_/a_219_297# 0.07fF
C5962 _349_/a_292_297# VPWR 0.01fF
C5963 _393_/A _631_/B 0.08fF
C5964 B[2] _610_/Y 0.17fF
C5965 _538_/A _559_/X 0.58fF
C5966 input7/a_27_47# _483_/X 0.02fF
C5967 _614_/a_76_199# _614_/a_226_297# 0.01fF
C5968 _614_/a_226_47# _614_/a_489_413# 0.02fF
C5969 _542_/A _486_/A 0.06fF
C5970 _396_/a_250_297# VPWR 0.75fF
C5971 _633_/Y B[7] 0.05fF
C5972 _446_/X _472_/Y 0.24fF
C5973 _585_/B _486_/X 1.26fF
C5974 _355_/A _346_/A 0.04fF
C5975 _485_/a_27_47# _547_/a_222_93# 0.00fF
C5976 _355_/A _478_/A 1.26fF
C5977 _469_/a_381_47# _610_/A 0.10fF
C5978 _613_/a_323_297# _433_/Y 0.03fF
C5979 _433_/Y _469_/X 2.62fF
C5980 _390_/D _542_/A 0.05fF
C5981 _576_/X _485_/D 0.35fF
C5982 _340_/A _390_/B 0.04fF
C5983 _557_/Y _582_/Y 0.43fF
C5984 _483_/a_93_21# _483_/a_250_297# 0.50fF
C5985 _411_/B _390_/D 0.05fF
C5986 _445_/X _390_/a_27_47# 0.05fF
C5987 _582_/Y _602_/A 1.34fF
C5988 _586_/S _469_/X 0.11fF
C5989 _487_/X _449_/A 0.49fF
C5990 input3/a_558_47# _390_/D 0.11fF
C5991 _599_/Y _624_/X 0.11fF
C5992 _524_/X _489_/X 0.02fF
C5993 input5/a_381_47# _390_/B 0.12fF
C5994 _454_/a_76_199# _454_/X 0.30fF
C5995 _494_/a_489_413# _492_/X 0.07fF
C5996 _453_/X _447_/B 0.00fF
C5997 _402_/a_27_47# _472_/B 0.30fF
C5998 _554_/B _556_/A 0.03fF
C5999 _379_/a_78_199# _448_/B 0.12fF
C6000 _545_/Y _572_/A 0.03fF
C6001 _391_/B _410_/C 0.09fF
C6002 _344_/a_78_199# _343_/X 0.30fF
C6003 _360_/a_76_199# _360_/a_226_47# 0.49fF
C6004 _446_/X _446_/a_250_297# 0.03fF
C6005 _626_/Y _468_/X 0.21fF
C6006 _368_/B _475_/A 0.01fF
C6007 _386_/a_558_47# _386_/a_841_47# 0.07fF
C6008 input7/a_27_47# A[6] 0.44fF
C6009 _363_/A _426_/A 0.09fF
C6010 _584_/a_150_297# _622_/X 0.01fF
C6011 _458_/a_78_199# VPWR 0.58fF
C6012 _594_/a_109_297# VPWR 0.39fF
C6013 _411_/A _409_/a_78_199# 0.21fF
C6014 _326_/A _409_/a_493_297# 0.08fF
C6015 _417_/a_27_47# _418_/B 0.18fF
C6016 _573_/A _595_/X 0.42fF
C6017 _583_/X input12/a_841_47# 0.05fF
C6018 _400_/a_80_21# _631_/B 0.11fF
C6019 output30/a_27_47# M[7] 0.48fF
C6020 _540_/X _469_/X 0.07fF
C6021 _594_/a_373_47# _573_/Y 0.02fF
C6022 _328_/X _329_/X 0.01fF
C6023 _519_/a_29_53# _519_/C 0.30fF
C6024 _475_/X _475_/a_68_297# 0.47fF
C6025 _417_/D _519_/C 0.00fF
C6026 _530_/a_556_47# _531_/B 0.02fF
C6027 _381_/C _449_/A 1.00fF
C6028 _461_/a_78_199# _461_/a_215_47# 0.26fF
C6029 _375_/a_448_47# _417_/A 0.02fF
C6030 _633_/a_74_47# _368_/B 0.31fF
C6031 _338_/a_544_297# VPWR 0.01fF
C6032 _360_/X _475_/A 0.75fF
C6033 _587_/A _533_/a_227_47# 0.02fF
C6034 _359_/X _454_/X 0.42fF
C6035 _614_/a_226_297# _611_/X 0.04fF
C6036 _614_/a_489_413# _613_/X 0.14fF
C6037 _386_/X _483_/a_250_297# 0.03fF
C6038 _563_/D _394_/a_381_47# 0.02fF
C6039 _544_/A _584_/A 1.68fF
C6040 _487_/X _517_/a_150_297# 0.03fF
C6041 _590_/A _590_/a_68_297# 0.36fF
C6042 _391_/A _442_/B 0.03fF
C6043 _600_/a_114_47# VPWR 0.01fF
C6044 _376_/X _420_/a_448_47# 0.14fF
C6045 _480_/A VPWR 1.03fF
C6046 _396_/X VPWR 1.04fF
C6047 _587_/a_27_47# _624_/a_76_199# 0.02fF
C6048 _513_/A _447_/X 0.25fF
C6049 _597_/a_78_199# _559_/X 0.59fF
C6050 _626_/Y _631_/Y 0.03fF
C6051 _470_/a_80_21# _470_/a_209_297# 0.16fF
C6052 _595_/a_77_199# _588_/A 0.45fF
C6053 _417_/D _539_/X 0.52fF
C6054 M[4] _432_/X 0.14fF
C6055 _533_/a_539_297# VPWR 0.02fF
C6056 _445_/X _446_/a_93_21# 0.21fF
C6057 _357_/a_27_47# _381_/B 0.41fF
C6058 _412_/a_226_47# _419_/X 0.02fF
C6059 _568_/a_323_297# _566_/Y 0.03fF
C6060 _445_/X _391_/B 0.21fF
C6061 _627_/C _564_/A 0.07fF
C6062 _386_/A _390_/a_27_47# 0.10fF
C6063 _503_/a_841_47# VPWR 0.43fF
C6064 _563_/A _547_/X 0.03fF
C6065 _517_/a_68_297# _380_/A 0.03fF
C6066 _454_/X _447_/X 0.50fF
C6067 _582_/Y _606_/A 0.43fF
C6068 _584_/A _391_/B 0.14fF
C6069 _438_/a_68_297# _438_/a_150_297# 0.02fF
C6070 VPWR _481_/A 7.22fF
C6071 _509_/Y _507_/Y 0.04fF
C6072 _360_/a_226_47# _353_/X 0.25fF
C6073 _433_/Y _546_/X 0.02fF
C6074 _447_/B _542_/D 1.59fF
C6075 _396_/a_93_21# _383_/X 0.01fF
C6076 _633_/Y VPWR 17.88fF
C6077 _631_/B _433_/Y 0.03fF
C6078 _408_/B _350_/C 1.08fF
C6079 _404_/a_62_47# _404_/a_381_47# 0.08fF
C6080 _627_/A _547_/X 0.03fF
C6081 _382_/X _383_/a_76_199# 0.24fF
C6082 _468_/X _527_/A 0.21fF
C6083 _439_/X _436_/a_68_297# 0.00fF
C6084 input15/a_75_212# B[6] 0.43fF
C6085 _337_/a_68_297# _337_/X 0.27fF
C6086 _563_/B _454_/X 1.36fF
C6087 _383_/a_226_47# _452_/A 0.06fF
C6088 _492_/a_226_47# _504_/X 0.06fF
C6089 _426_/A _374_/X 0.26fF
C6090 _544_/A _386_/A 0.06fF
C6091 _378_/A _512_/a_78_199# 0.01fF
C6092 _426_/a_68_297# _426_/a_150_297# 0.02fF
C6093 _375_/X _359_/A 0.20fF
C6094 _490_/a_215_47# VPWR 0.14fF
C6095 _540_/X _546_/X 0.03fF
C6096 _548_/X _547_/X 0.64fF
C6097 _518_/a_250_297# _515_/A 0.10fF
C6098 _408_/B _367_/C 0.80fF
C6099 _613_/X _503_/A 0.02fF
C6100 _330_/A _442_/B 0.70fF
C6101 _576_/X _598_/B 0.13fF
C6102 _630_/a_76_199# _630_/a_489_413# 0.12fF
C6103 _617_/a_113_297# _616_/B 0.09fF
C6104 _617_/a_199_47# _616_/A 0.14fF
C6105 _575_/X _574_/X 1.71fF
C6106 _350_/C _445_/a_68_297# 0.00fF
C6107 _487_/X _417_/D 2.29fF
C6108 _509_/Y _511_/a_256_47# 0.03fF
C6109 _362_/a_226_47# _362_/a_489_413# 0.02fF
C6110 _362_/a_76_199# _362_/a_226_297# 0.01fF
C6111 _519_/X _486_/A 0.22fF
C6112 _510_/A _436_/X 0.03fF
C6113 _386_/A _446_/a_93_21# 0.01fF
C6114 _451_/A _563_/B 0.02fF
C6115 _562_/a_78_199# _563_/A 0.01fF
C6116 A[4] _478_/A 0.06fF
C6117 _487_/X _347_/A 0.52fF
C6118 _475_/X _468_/a_78_199# 0.01fF
C6119 _491_/X _489_/X 0.82fF
C6120 _533_/X _454_/X 0.36fF
C6121 _534_/a_80_21# _386_/a_62_47# 0.02fF
C6122 _554_/A _555_/a_27_413# 0.22fF
C6123 _460_/a_489_413# VPWR 0.39fF
C6124 _386_/A _391_/B 0.19fF
C6125 _503_/A _609_/a_80_21# 0.16fF
C6126 _629_/A _371_/A 0.02fF
C6127 _417_/A _351_/A 0.07fF
C6128 _554_/X _554_/B 0.60fF
C6129 _464_/A _464_/Y 0.59fF
C6130 _579_/X _581_/B 1.40fF
C6131 _488_/a_76_199# _627_/A 0.08fF
C6132 _441_/a_493_297# _340_/A 0.01fF
C6133 _519_/a_29_53# _519_/a_183_297# 0.04fF
C6134 _426_/a_68_297# _427_/A 0.27fF
C6135 _360_/X _390_/B 0.26fF
C6136 _442_/A _472_/B 0.44fF
C6137 _519_/a_29_53# _381_/C 0.04fF
C6138 _444_/A _410_/C 0.59fF
C6139 _410_/a_27_47# _631_/Y 0.22fF
C6140 _626_/Y _624_/a_489_47# 0.09fF
C6141 _561_/A _454_/a_76_199# 0.01fF
C6142 _533_/a_77_199# _533_/a_227_297# 0.13fF
C6143 _476_/X _446_/X 0.03fF
C6144 _368_/a_68_297# _368_/A 0.45fF
C6145 _417_/D _381_/C 0.04fF
C6146 _411_/B _411_/a_68_297# 0.36fF
C6147 _625_/a_277_47# _601_/A 0.09fF
C6148 _426_/B _466_/X 0.35fF
C6149 _430_/A VPWR 1.74fF
C6150 _609_/a_80_21# _609_/a_209_297# 0.16fF
C6151 _611_/a_27_297# _627_/C 0.37fF
C6152 _633_/A _631_/A 0.01fF
C6153 _375_/X _367_/C 0.53fF
C6154 _390_/B _465_/X 0.06fF
C6155 B[7] _454_/a_76_199# 0.07fF
C6156 _347_/a_27_47# _378_/A 0.16fF
C6157 _536_/Y _390_/D 0.05fF
C6158 _616_/B _601_/A 0.25fF
C6159 _616_/A _624_/X 0.07fF
C6160 _587_/A _599_/Y 0.39fF
C6161 _463_/a_226_47# _497_/A 0.01fF
C6162 _615_/a_493_297# VPWR 0.02fF
C6163 B[7] _585_/B 0.08fF
C6164 B[1] _335_/a_841_47# 0.09fF
C6165 _454_/X _322_/a_27_47# 0.10fF
C6166 _436_/A _458_/X 0.42fF
C6167 _510_/a_68_297# VPWR 0.31fF
C6168 _421_/a_556_47# _631_/B 0.02fF
C6169 VPWR _413_/a_68_297# 0.28fF
C6170 _417_/D _570_/A 0.23fF
C6171 _544_/A _386_/X 0.00fF
C6172 _324_/a_558_47# _324_/a_664_47# 0.60fF
C6173 _324_/a_381_47# _324_/a_841_47# 0.03fF
C6174 _590_/B _588_/Y 0.21fF
C6175 _516_/A _356_/a_78_199# 0.34fF
C6176 _445_/A _409_/a_493_297# 0.02fF
C6177 _474_/A _510_/A 0.24fF
C6178 _550_/X _511_/X 0.03fF
C6179 _356_/a_493_297# _481_/A 0.08fF
C6180 _567_/Y _587_/A 0.44fF
C6181 _524_/X _554_/a_68_297# 0.01fF
C6182 _347_/A _570_/A 0.05fF
C6183 _542_/C _417_/D 0.10fF
C6184 _418_/a_68_297# _418_/X 0.33fF
C6185 _611_/a_27_297# _611_/a_109_297# 0.45fF
C6186 _542_/A _628_/Y 0.03fF
C6187 _403_/a_27_47# _539_/A 0.07fF
C6188 _578_/a_493_297# _550_/X 0.08fF
C6189 _578_/a_78_199# _580_/B 0.21fF
C6190 _578_/a_215_47# _551_/X 0.18fF
C6191 _374_/a_78_199# _374_/a_215_47# 0.26fF
C6192 B[0] _587_/A 0.05fF
C6193 _360_/X _328_/B 1.14fF
C6194 _444_/A _445_/X 0.18fF
C6195 _380_/A _408_/B 0.03fF
C6196 _469_/a_664_47# _586_/a_505_21# 0.01fF
C6197 _386_/X _446_/a_93_21# 0.46fF
C6198 _580_/B _606_/A 1.27fF
C6199 _543_/Y VPWR 0.50fF
C6200 _616_/A _622_/C 0.00fF
C6201 _623_/X _588_/A 0.60fF
C6202 _454_/X _509_/Y 0.41fF
C6203 _369_/a_76_199# _329_/X 0.01fF
C6204 _369_/a_489_413# _343_/X 0.14fF
C6205 _544_/a_381_47# _588_/A 0.61fF
C6206 _515_/Y VPWR 0.84fF
C6207 _532_/a_76_199# _528_/a_299_297# 0.02fF
C6208 _532_/a_206_369# _528_/a_81_21# 0.01fF
C6209 _456_/a_76_199# _456_/a_226_297# 0.01fF
C6210 _456_/a_226_47# _456_/a_489_413# 0.02fF
C6211 _386_/X _391_/B 0.72fF
C6212 VPWR _602_/Y 1.37fF
C6213 _627_/C _454_/X 0.03fF
C6214 _561_/A _447_/X 0.05fF
C6215 _587_/A _468_/a_493_297# 0.02fF
C6216 _563_/B _627_/B 0.05fF
C6217 _567_/B _469_/A 0.08fF
C6218 _595_/a_77_199# _571_/a_93_21# 0.02fF
C6219 _424_/a_76_199# _424_/a_226_47# 0.49fF
C6220 _335_/a_664_47# _417_/A 0.20fF
C6221 _448_/A _448_/B 0.19fF
C6222 _390_/B M[10] 0.28fF
C6223 _542_/D _486_/B 0.02fF
C6224 _583_/X M[1] 0.05fF
C6225 _620_/X _616_/Y 1.29fF
C6226 _452_/X _542_/A 0.19fF
C6227 B[7] _447_/X 0.63fF
C6228 VPWR _521_/a_78_199# 0.63fF
C6229 _542_/B _442_/B 0.36fF
C6230 _476_/X _492_/a_76_199# 0.33fF
C6231 _628_/a_734_297# _628_/a_300_47# 0.03fF
C6232 _626_/a_109_47# _623_/X 0.23fF
C6233 input6/a_27_47# _380_/A 0.22fF
C6234 _520_/a_226_47# _381_/B 0.14fF
C6235 _476_/a_346_47# _390_/B 0.02fF
C6236 _436_/A _395_/a_68_297# 0.42fF
C6237 _549_/X _549_/a_226_47# 0.05fF
C6238 VPWR _468_/a_292_297# 0.01fF
C6239 _622_/a_29_53# _622_/C 0.30fF
C6240 _343_/a_226_47# _338_/X 0.61fF
C6241 _584_/A _394_/a_558_47# 0.11fF
C6242 _418_/X _542_/D 0.06fF
C6243 _458_/X _478_/A 0.03fF
C6244 _436_/A _350_/B 2.13fF
C6245 _462_/X _460_/X 0.08fF
C6246 _627_/C _451_/A 0.30fF
C6247 _497_/A _498_/A 0.67fF
C6248 _561_/A _563_/B 0.36fF
C6249 _569_/Y _469_/X 0.92fF
C6250 _375_/X _380_/A 0.03fF
C6251 B[7] _616_/Y 0.20fF
C6252 _520_/X _515_/A 0.91fF
C6253 _433_/Y output29/a_27_47# 0.43fF
C6254 _379_/a_215_47# _356_/a_215_47# 0.02fF
C6255 _630_/a_76_199# _629_/a_68_297# 0.02fF
C6256 _419_/X _332_/X 0.03fF
C6257 _563_/B B[7] 1.22fF
C6258 _338_/a_79_199# _366_/a_76_199# 0.03fF
C6259 _482_/X _410_/C 0.42fF
C6260 _605_/a_80_21# _582_/Y 0.02fF
C6261 _582_/a_109_297# VPWR 0.01fF
C6262 _417_/A _519_/A 3.46fF
C6263 _542_/D _622_/C 0.09fF
C6264 _352_/X _371_/B 0.03fF
C6265 _431_/a_76_199# _390_/B 0.10fF
C6266 _454_/a_76_199# VPWR 0.58fF
C6267 _444_/A _386_/A 0.21fF
C6268 _387_/a_78_199# _584_/A 0.08fF
C6269 _410_/B _446_/a_93_21# 0.42fF
C6270 _448_/a_68_297# _542_/D 0.20fF
C6271 _520_/X _535_/Y 0.48fF
C6272 VPWR _558_/a_227_297# 0.01fF
C6273 _627_/a_27_297# _627_/a_277_297# 0.05fF
C6274 _620_/a_76_199# _620_/X 0.22fF
C6275 _620_/a_226_47# _618_/Y 0.31fF
C6276 _368_/a_68_297# _370_/A 0.27fF
C6277 _455_/a_79_199# _455_/a_222_93# 0.51fF
C6278 _585_/B VPWR 5.05fF
C6279 _442_/D _546_/a_489_413# 0.09fF
C6280 _375_/X _384_/a_226_47# 0.22fF
C6281 _540_/a_346_47# _469_/X 0.03fF
C6282 _613_/a_227_47# _627_/D 0.11fF
C6283 _493_/a_215_47# _457_/X 0.11fF
C6284 _590_/a_68_297# _590_/a_150_297# 0.02fF
C6285 _566_/A _571_/a_584_47# 0.02fF
C6286 _487_/X _477_/a_78_199# 0.12fF
C6287 _459_/a_76_199# _460_/a_226_47# 0.01fF
C6288 _459_/a_226_47# _460_/a_76_199# 0.01fF
C6289 B[1] _363_/A 0.33fF
C6290 _505_/a_80_21# _505_/a_303_47# 0.04fF
C6291 _375_/a_222_93# _375_/X 0.06fF
C6292 _591_/Y _613_/X 0.05fF
C6293 _352_/X _361_/a_489_413# 0.07fF
C6294 B[1] _420_/X 0.08fF
C6295 _469_/a_558_47# _586_/a_76_199# 0.00fF
C6296 _583_/X _622_/X 0.01fF
C6297 _527_/B _531_/B 0.12fF
C6298 _350_/B _350_/X 0.02fF
C6299 M[7] _557_/B 1.15fF
C6300 _363_/a_68_297# _363_/B 0.33fF
C6301 _510_/A _385_/a_558_47# 0.07fF
C6302 _359_/X VPWR 1.73fF
C6303 _611_/X _590_/B 0.20fF
C6304 _386_/A _394_/a_558_47# 0.01fF
C6305 _563_/A _481_/A 1.89fF
C6306 _351_/A _631_/B 0.09fF
C6307 _338_/a_79_199# _631_/B 0.06fF
C6308 _386_/a_841_47# VPWR 0.33fF
C6309 _572_/B _574_/a_81_21# 0.02fF
C6310 _337_/B _367_/C 0.01fF
C6311 _563_/A _633_/Y 0.04fF
C6312 _350_/a_27_297# _313_/A 0.01fF
C6313 _422_/a_226_47# _421_/a_76_199# 0.01fF
C6314 _566_/A _546_/a_226_297# 0.01fF
C6315 _607_/X _612_/Y 0.03fF
C6316 _448_/A _453_/a_93_21# 0.04fF
C6317 _608_/X _627_/B 0.01fF
C6318 _537_/a_77_199# _537_/a_323_297# 0.05fF
C6319 _476_/a_93_21# _475_/X 0.21fF
C6320 _390_/D _539_/A 0.03fF
C6321 _455_/X _472_/B 0.03fF
C6322 _347_/A _477_/a_493_297# 0.08fF
C6323 _563_/D _442_/B 0.12fF
C6324 _365_/a_81_21# _363_/B 0.02fF
C6325 _493_/a_78_199# _458_/X 0.27fF
C6326 _493_/a_215_47# _459_/X 0.05fF
C6327 _519_/A _484_/a_215_47# 0.05fF
C6328 _425_/a_489_413# _424_/X 0.14fF
C6329 _627_/A _633_/Y 0.27fF
C6330 _410_/C _539_/X 0.14fF
C6331 _509_/A _472_/B 0.29fF
C6332 _627_/C _627_/B 1.39fF
C6333 _447_/X VPWR 1.95fF
C6334 _583_/X _580_/a_68_297# 0.20fF
C6335 _334_/a_197_47# VPWR 0.02fF
C6336 M[2] _338_/X 0.44fF
C6337 _569_/Y _546_/X 0.09fF
C6338 _420_/X _383_/X 0.03fF
C6339 _612_/A _616_/A 0.26fF
C6340 _360_/X _361_/a_226_47# 0.56fF
C6341 VPWR _625_/a_27_297# 1.44fF
C6342 _556_/Y M[7] 0.20fF
C6343 _599_/A _597_/a_215_47# 0.03fF
C6344 _391_/B _395_/X 0.16fF
C6345 _365_/a_384_47# _432_/B 0.02fF
C6346 _328_/A _328_/a_68_297# 0.33fF
C6347 VPWR _558_/X 3.63fF
C6348 _618_/Y _619_/Y 1.33fF
C6349 output17/a_27_47# _552_/a_76_199# 0.01fF
C6350 _375_/X _455_/X 0.38fF
C6351 _469_/a_62_47# _545_/Y 0.14fF
C6352 _347_/A _518_/a_256_47# 0.03fF
C6353 _464_/A _500_/a_215_47# 0.10fF
C6354 _444_/A _386_/X 0.06fF
C6355 _423_/X VPWR 3.98fF
C6356 _385_/a_381_47# _475_/A 0.12fF
C6357 _625_/Y _625_/a_27_47# 0.03fF
C6358 _553_/a_215_47# _524_/X 0.10fF
C6359 _587_/A _572_/A 0.47fF
C6360 _544_/A M[9] 0.47fF
C6361 _417_/D _540_/a_93_21# 0.21fF
C6362 _494_/a_489_413# _626_/Y 0.09fF
C6363 VPWR _409_/a_292_297# 0.01fF
C6364 VPWR _616_/Y 3.35fF
C6365 M[13] _442_/D 0.10fF
C6366 _408_/X _393_/A 0.03fF
C6367 _381_/C _547_/a_79_199# 0.17fF
C6368 _567_/B _459_/a_76_199# 0.08fF
C6369 input5/a_664_47# _430_/X 0.01fF
C6370 input5/a_558_47# _428_/X 0.00fF
C6371 _349_/a_78_199# _349_/a_292_297# 0.03fF
C6372 _561_/A _627_/C 0.02fF
C6373 _563_/B VPWR 6.47fF
C6374 _573_/Y _616_/B 0.00fF
C6375 _392_/A _631_/A 0.10fF
C6376 _623_/X _616_/B 0.14fF
C6377 _625_/Y _616_/A 0.66fF
C6378 _336_/a_292_297# _442_/B 0.02fF
C6379 _398_/a_226_47# _399_/a_78_199# 0.01fF
C6380 _518_/a_93_21# _570_/A 0.03fF
C6381 _627_/C B[7] 1.36fF
C6382 _436_/A _587_/A 0.40fF
C6383 _627_/A _475_/a_150_297# 0.02fF
C6384 _572_/B VPWR 1.66fF
C6385 _396_/a_93_21# _396_/a_250_297# 0.50fF
C6386 _386_/a_381_47# _381_/B 0.01fF
C6387 M[8] _466_/X 0.52fF
C6388 _408_/B _336_/a_215_47# 0.07fF
C6389 _507_/Y _469_/X 0.09fF
C6390 _612_/A _620_/a_226_47# 0.08fF
C6391 _386_/A _482_/X 0.10fF
C6392 _352_/X _361_/a_76_199# 0.32fF
C6393 VPWR _550_/a_78_199# 0.62fF
C6394 _625_/Y _572_/A 0.17fF
C6395 _416_/a_78_199# _416_/a_292_297# 0.03fF
C6396 _416_/a_215_47# _448_/B 0.13fF
C6397 _327_/a_215_47# VPWR 0.04fF
C6398 _623_/a_76_199# _621_/X 0.46fF
C6399 _461_/a_215_47# _461_/X 0.01fF
C6400 _501_/Y _558_/X 0.05fF
C6401 _487_/X _410_/C 0.13fF
C6402 _503_/A _571_/a_250_297# 0.14fF
C6403 _533_/X VPWR 4.22fF
C6404 _626_/Y _522_/X 0.42fF
C6405 _520_/X A[3] 0.47fF
C6406 _313_/A _475_/A 0.72fF
C6407 _620_/a_76_199# VPWR 0.47fF
C6408 _590_/A A[3] 0.09fF
C6409 _611_/a_109_297# B[7] 0.06fF
C6410 _375_/X _397_/a_76_199# 0.01fF
C6411 _382_/X _420_/a_222_93# 0.11fF
C6412 _380_/A _517_/X 0.11fF
C6413 _567_/B _502_/a_78_199# 0.18fF
C6414 _474_/A _472_/Y 1.19fF
C6415 _485_/a_27_47# _485_/a_109_47# 0.03fF
C6416 _543_/B _512_/a_78_199# 0.01fF
C6417 _411_/B _437_/a_448_47# 0.08fF
C6418 _513_/A _417_/A 0.57fF
C6419 _628_/a_300_47# VPWR 0.08fF
C6420 _444_/A _410_/B 1.69fF
C6421 _441_/a_215_47# _346_/A 0.10fF
C6422 _442_/D _442_/A 0.49fF
C6423 _417_/a_27_47# _367_/C 0.10fF
C6424 _482_/X _483_/a_93_21# 0.21fF
C6425 _381_/C _410_/C 0.64fF
C6426 _538_/Y _469_/X 0.36fF
C6427 _476_/a_250_297# VPWR 0.74fF
C6428 _511_/a_256_47# _469_/X 0.04fF
C6429 _540_/a_250_297# _472_/B 0.09fF
C6430 _461_/a_215_47# _407_/a_27_47# 0.06fF
C6431 _371_/B _350_/X 0.41fF
C6432 _436_/X _437_/X 0.03fF
C6433 _519_/A _631_/B 0.02fF
C6434 _328_/B _314_/a_68_297# 0.01fF
C6435 _542_/D _514_/a_68_297# 0.02fF
C6436 _542_/A _447_/B 0.40fF
C6437 _623_/a_76_199# _623_/a_226_47# 0.49fF
C6438 _417_/A _454_/X 0.15fF
C6439 _587_/A _478_/A 0.50fF
C6440 _425_/a_76_199# _478_/A 0.08fF
C6441 _503_/A _535_/Y 0.73fF
C6442 VPWR _322_/a_27_47# 0.70fF
C6443 VPWR _553_/a_292_297# 0.01fF
C6444 _452_/a_150_297# _628_/Y 0.01fF
C6445 _429_/a_76_199# _429_/a_489_413# 0.12fF
C6446 _330_/A _384_/a_489_413# 0.02fF
C6447 _612_/Y _588_/A 0.39fF
C6448 _396_/a_93_21# _396_/X 0.19fF
C6449 _392_/A _391_/a_68_297# 0.27fF
C6450 _499_/a_299_297# _498_/Y 0.07fF
C6451 _567_/Y _433_/Y 0.21fF
C6452 input3/a_841_47# _485_/D 0.05fF
C6453 _390_/D _588_/A 0.26fF
C6454 _595_/a_227_47# VPWR 0.04fF
C6455 _475_/X _504_/a_539_297# 0.03fF
C6456 _543_/Y _627_/A 0.11fF
C6457 _612_/A _619_/Y 0.50fF
C6458 _410_/C _570_/A 0.00fF
C6459 B[0] _433_/Y 0.08fF
C6460 _594_/a_27_297# _594_/a_109_297# 0.45fF
C6461 _422_/a_76_199# _422_/a_489_413# 0.12fF
C6462 _487_/X _584_/A 0.69fF
C6463 _537_/a_323_297# VPWR 0.02fF
C6464 _545_/a_109_297# _610_/A 0.01fF
C6465 _404_/a_381_47# _543_/A 0.07fF
C6466 _410_/C _316_/a_62_47# 0.31fF
C6467 _583_/X _599_/A 0.03fF
C6468 _608_/X VPWR 1.01fF
C6469 _542_/C _410_/C 1.15fF
C6470 _386_/X _482_/X 0.07fF
C6471 VPWR _369_/a_226_47# 0.06fF
C6472 _358_/a_27_47# _359_/A 0.01fF
C6473 _375_/X _335_/a_381_47# 0.16fF
C6474 A[6] _449_/A 0.03fF
C6475 _509_/Y VPWR 1.28fF
C6476 B[6] _531_/B 0.08fF
C6477 _370_/a_68_297# VPWR 0.25fF
C6478 _567_/B _547_/X 0.06fF
C6479 _567_/Y _540_/X 0.20fF
C6480 _469_/X _486_/X 0.09fF
C6481 _519_/X _520_/a_226_47# 0.69fF
C6482 _525_/a_76_199# _525_/a_489_413# 0.12fF
C6483 _392_/Y _631_/A 0.01fF
C6484 _490_/X _456_/X 0.10fF
C6485 _627_/C VPWR 6.80fF
C6486 _468_/a_215_47# VPWR 0.05fF
C6487 _381_/B _486_/B 0.10fF
C6488 _381_/C _584_/A 0.47fF
C6489 _357_/a_27_47# _539_/A 0.01fF
C6490 B[0] _540_/X 0.05fF
C6491 _527_/Y _527_/a_109_297# 0.02fF
C6492 _487_/a_215_47# _454_/a_76_199# 0.01fF
C6493 _601_/Y _619_/Y 0.03fF
C6494 _426_/B _431_/X 0.01fF
C6495 _373_/a_113_297# _371_/A 0.13fF
C6496 _338_/a_79_199# _338_/a_448_47# 0.13fF
C6497 _610_/A _588_/Y 0.10fF
C6498 _544_/A _515_/A 0.08fF
C6499 _411_/A _470_/a_209_297# 0.13fF
C6500 _424_/X _407_/Y 1.56fF
C6501 _483_/a_584_47# _542_/A 0.04fF
C6502 _604_/a_80_21# _557_/B 0.31fF
C6503 _469_/a_664_47# _503_/A 0.06fF
C6504 _347_/A _510_/A 0.16fF
C6505 _350_/a_27_297# _408_/B 0.15fF
C6506 _417_/A _337_/A 0.03fF
C6507 _454_/X _469_/X 0.08fF
C6508 _510_/A _332_/X 0.20fF
C6509 _611_/a_109_297# VPWR 0.39fF
C6510 _313_/A _390_/B 0.34fF
C6511 _582_/Y _556_/A 0.05fF
C6512 _472_/a_109_297# VPWR 0.01fF
C6513 _584_/A _570_/A 0.22fF
C6514 _436_/A _393_/A 0.03fF
C6515 _519_/a_29_53# _485_/D 0.02fF
C6516 _534_/a_303_47# _515_/A 0.01fF
C6517 _542_/C _445_/X 0.53fF
C6518 _429_/a_489_413# VPWR 0.39fF
C6519 _417_/D _485_/D 0.12fF
C6520 _542_/B _520_/X 0.03fF
C6521 _487_/X _386_/A 0.14fF
C6522 _627_/A _585_/B 0.75fF
C6523 _488_/a_226_47# _507_/Y 0.01fF
C6524 _458_/a_215_47# _421_/X 0.05fF
C6525 _455_/X _446_/X 0.09fF
C6526 _459_/a_489_413# _458_/X 0.14fF
C6527 _518_/a_93_21# _518_/a_256_47# 0.03fF
C6528 _347_/A _485_/D 0.03fF
C6529 _404_/a_62_47# _585_/B 0.62fF
C6530 _479_/B _505_/a_80_21# 0.40fF
C6531 _358_/a_27_47# _442_/A 0.29fF
C6532 _631_/Y _539_/A 0.05fF
C6533 _359_/B _359_/A 1.25fF
C6534 _487_/X _521_/X 0.01fF
C6535 _629_/A _365_/a_81_21# 0.48fF
C6536 _423_/a_292_297# _384_/X 0.02fF
C6537 _556_/Y _604_/a_80_21# 0.28fF
C6538 _417_/D _483_/X 0.29fF
C6539 _631_/Y _489_/X 0.03fF
C6540 _598_/B _593_/Y 0.26fF
C6541 _359_/a_68_297# _381_/C 0.00fF
C6542 _504_/a_227_47# VPWR 0.04fF
C6543 _362_/a_76_199# _352_/X 0.01fF
C6544 _342_/X _369_/a_226_47# 0.40fF
C6545 _478_/A _466_/a_78_199# 0.17fF
C6546 _487_/a_215_47# _447_/X 0.33fF
C6547 _503_/a_664_47# _503_/a_841_47# 0.29fF
C6548 _501_/a_109_47# _501_/a_397_297# 0.05fF
C6549 _503_/A A[3] 2.47fF
C6550 B[2] _620_/X 0.07fF
C6551 _390_/D _559_/X 3.09fF
C6552 _528_/a_299_297# _530_/X 0.03fF
C6553 _436_/A _400_/a_80_21# 0.00fF
C6554 _524_/a_78_199# VPWR 0.57fF
C6555 _538_/A _472_/B 0.11fF
C6556 _448_/B _356_/a_78_199# 0.01fF
C6557 _516_/a_27_47# _481_/A 0.01fF
C6558 _631_/A _332_/X 0.67fF
C6559 _425_/a_226_297# VPWR 0.00fF
C6560 _542_/D _484_/a_78_199# 0.01fF
C6561 _481_/a_27_47# _539_/A 0.29fF
C6562 _336_/a_215_47# _337_/B 0.01fF
C6563 _386_/A _570_/A 0.44fF
C6564 VPWR _501_/a_397_297# 0.53fF
C6565 _542_/A _486_/B 0.14fF
C6566 _584_/A _419_/X 0.32fF
C6567 _474_/A _476_/X 0.06fF
C6568 _570_/B _587_/A 0.50fF
C6569 _422_/X _433_/Y 0.15fF
C6570 _626_/Y _587_/A 0.04fF
C6571 _612_/Y _625_/a_277_47# 0.02fF
C6572 _419_/X _420_/a_79_199# 0.17fF
C6573 _384_/X input14/a_27_47# 0.01fF
C6574 _487_/a_215_47# _563_/B 0.12fF
C6575 _574_/X _575_/a_493_297# 0.02fF
C6576 _542_/C _386_/A 2.13fF
C6577 _575_/X _575_/a_215_47# 0.01fF
C6578 _607_/X _607_/a_215_47# 0.01fF
C6579 _417_/D A[6] 0.03fF
C6580 _626_/Y _612_/A 0.09fF
C6581 _563_/A _563_/B 0.82fF
C6582 _455_/X _442_/D 1.14fF
C6583 _557_/A VPWR 3.78fF
C6584 _605_/a_209_297# _604_/X 0.06fF
C6585 _544_/A _447_/a_68_297# 0.34fF
C6586 _352_/X _374_/a_78_199# 0.01fF
C6587 _440_/a_226_47# _436_/X 0.25fF
C6588 _386_/X _487_/X 0.11fF
C6589 _408_/B _475_/A 0.42fF
C6590 _603_/Y _602_/Y 1.01fF
C6591 _518_/a_250_297# _518_/X 0.03fF
C6592 _347_/A A[6] 0.05fF
C6593 _612_/Y _616_/B 0.47fF
C6594 A[2] _618_/A 0.00fF
C6595 _503_/a_62_47# _446_/X 0.14fF
C6596 _513_/a_197_47# _542_/B 0.12fF
C6597 _359_/B _442_/A 0.08fF
C6598 _585_/B _537_/a_227_47# 0.01fF
C6599 _360_/X _332_/a_68_297# 0.20fF
C6600 _363_/A _432_/B 0.80fF
C6601 _524_/a_215_47# _476_/X 0.29fF
C6602 _493_/X _502_/a_215_47# 0.10fF
C6603 _478_/a_27_47# _478_/a_109_47# 0.03fF
C6604 _572_/A _433_/Y 0.02fF
C6605 _593_/A _622_/C 0.09fF
C6606 _391_/A _391_/B 0.17fF
C6607 _563_/D _520_/X 0.03fF
C6608 _611_/X _610_/A 0.41fF
C6609 _516_/A _355_/A 0.01fF
C6610 _518_/X _547_/a_222_93# 0.03fF
C6611 _625_/Y _626_/Y 0.29fF
C6612 _488_/a_226_47# _486_/X 0.31fF
C6613 _586_/S _572_/A 0.32fF
C6614 _374_/a_493_297# _374_/X 0.02fF
C6615 _475_/A _472_/B 0.20fF
C6616 _386_/A _535_/A 0.03fF
C6617 _544_/A _378_/a_558_47# 0.11fF
C6618 _490_/a_78_199# _489_/X 0.01fF
C6619 _335_/a_841_47# _633_/Y 0.07fF
C6620 _431_/a_226_47# _428_/X 0.25fF
C6621 _431_/a_489_413# _430_/X 0.14fF
C6622 _360_/X _328_/A 0.03fF
C6623 _406_/A _436_/X 0.00fF
C6624 _540_/a_93_21# _410_/C 0.29fF
C6625 _501_/a_397_297# _501_/Y 0.26fF
C6626 _627_/B _469_/X 0.00fF
C6627 _544_/A _382_/B 0.02fF
C6628 _436_/A _433_/Y 0.03fF
C6629 _583_/X output23/a_27_47# 0.02fF
C6630 _475_/a_68_297# _633_/Y 0.01fF
C6631 _585_/B _508_/a_227_47# 0.11fF
C6632 _608_/a_78_199# _586_/S 0.12fF
C6633 _533_/X _627_/A 0.16fF
C6634 _485_/A _383_/X 0.70fF
C6635 _627_/A _473_/a_227_47# 0.02fF
C6636 _561_/A _484_/a_215_47# 0.03fF
C6637 _564_/a_219_297# _627_/D 0.00fF
C6638 _379_/a_215_47# _481_/A 0.01fF
C6639 _554_/X _582_/Y 0.36fF
C6640 _375_/X _475_/A 0.03fF
C6641 _587_/A _381_/B 0.10fF
C6642 _564_/a_27_53# _621_/X 0.02fF
C6643 _610_/A _618_/A 0.06fF
C6644 _610_/Y _616_/A 0.17fF
C6645 _586_/S _542_/D 0.79fF
C6646 _516_/A _520_/a_226_47# 0.04fF
C6647 _386_/X _570_/A 0.86fF
C6648 _439_/X _436_/X 1.58fF
C6649 _341_/a_27_47# _631_/B 0.22fF
C6650 _542_/C _386_/X 0.19fF
C6651 _476_/a_250_297# _627_/A 0.01fF
C6652 _569_/A _442_/D 0.02fF
C6653 B[7] _469_/X 0.01fF
C6654 _520_/X _518_/a_250_297# 0.26fF
C6655 _520_/a_76_199# _517_/X 0.05fF
C6656 _590_/A _586_/a_505_21# 0.14fF
C6657 _525_/a_489_413# _492_/a_226_47# 0.00fF
C6658 _420_/X _458_/a_78_199# 0.13fF
C6659 _337_/A _631_/B 0.80fF
C6660 _510_/A _336_/a_78_199# 0.13fF
C6661 _394_/a_381_47# _394_/a_558_47# 0.32fF
C6662 _322_/A _563_/D 0.03fF
C6663 _583_/X M[6] 0.49fF
C6664 _496_/a_292_297# _462_/X 0.08fF
C6665 _417_/D _418_/B 0.80fF
C6666 _330_/A _391_/B 0.47fF
C6667 _633_/A _367_/C 0.11fF
C6668 _496_/a_78_199# _461_/X 0.13fF
C6669 _460_/X _462_/a_489_413# 0.07fF
C6670 _561_/A _512_/a_78_199# 0.48fF
C6671 M[6] _622_/X 0.30fF
C6672 _475_/a_68_297# _475_/a_150_297# 0.02fF
C6673 _494_/X _492_/X 1.20fF
C6674 _533_/a_77_199# VPWR 0.95fF
C6675 _629_/X _426_/A 0.51fF
C6676 _410_/B _381_/C 0.66fF
C6677 _525_/X _554_/B 0.01fF
C6678 _527_/Y VPWR 1.93fF
C6679 _566_/Y A[3] 0.19fF
C6680 _469_/a_62_47# _587_/A 0.10fF
C6681 _432_/B _374_/X 0.01fF
C6682 input2/a_27_47# M[10] 0.10fF
C6683 _353_/X _375_/a_79_199# 0.03fF
C6684 _460_/a_226_47# _460_/a_489_413# 0.02fF
C6685 _460_/a_76_199# _460_/a_226_297# 0.01fF
C6686 _569_/A _588_/Y 0.02fF
C6687 _469_/a_62_47# _612_/A 0.01fF
C6688 _627_/A _595_/a_227_47# 0.11fF
C6689 VPWR _466_/a_215_47# 0.06fF
C6690 B[2] VPWR 2.34fF
C6691 _396_/X _363_/A 0.05fF
C6692 _433_/Y _478_/A 0.03fF
C6693 _584_/A _621_/X 0.23fF
C6694 _523_/a_489_413# _511_/X 0.07fF
C6695 _523_/a_226_47# _522_/X 0.50fF
C6696 _590_/A _591_/A 0.11fF
C6697 _417_/A VPWR 5.54fF
C6698 _506_/A _482_/X 0.24fF
C6699 _542_/a_27_47# _542_/D 0.25fF
C6700 _442_/D _627_/D 0.25fF
C6701 _516_/a_27_47# _515_/Y 0.01fF
C6702 _408_/B _390_/B 0.01fF
C6703 _563_/A _627_/C 2.10fF
C6704 _608_/X _627_/A 0.30fF
C6705 _530_/X _486_/A 0.08fF
C6706 _375_/a_222_93# _359_/B 0.06fF
C6707 _567_/B _633_/Y 1.43fF
C6708 _627_/A _509_/Y 0.10fF
C6709 _386_/X _419_/X 0.76fF
C6710 _390_/D _530_/X 0.03fF
C6711 output21/a_27_47# _625_/Y 0.01fF
C6712 _425_/a_489_413# _407_/Y 0.04fF
C6713 _546_/a_226_47# _515_/A 0.01fF
C6714 _473_/a_77_199# _472_/B 0.34fF
C6715 _627_/C _627_/A 1.17fF
C6716 _340_/A _355_/A 0.49fF
C6717 _410_/B _316_/a_62_47# 0.16fF
C6718 _385_/a_558_47# _394_/a_664_47# 0.01fF
C6719 _433_/a_109_47# _433_/Y 0.47fF
C6720 _519_/X _486_/B 0.17fF
C6721 _390_/a_27_47# _442_/B 0.02fF
C6722 _390_/B _472_/B 0.44fF
C6723 _351_/a_219_297# _350_/X 0.02fF
C6724 _410_/B _542_/C 0.23fF
C6725 _542_/B _390_/a_27_47# 0.39fF
C6726 _627_/D _588_/Y 1.63fF
C6727 _378_/A _542_/D 0.99fF
C6728 _412_/X VPWR 1.51fF
C6729 _546_/a_76_199# _546_/a_226_47# 0.49fF
C6730 _371_/a_68_297# _371_/a_150_297# 0.02fF
C6731 _336_/a_78_199# _631_/A 0.01fF
C6732 _633_/Y _420_/X 0.03fF
C6733 _587_/A _593_/A 0.23fF
C6734 _520_/X _518_/X 0.41fF
C6735 _417_/A _314_/X 0.51fF
C6736 _315_/a_161_47# B[7] 0.17fF
C6737 B[0] _540_/a_346_47# 0.02fF
C6738 _587_/A _542_/A 0.50fF
C6739 _567_/B _490_/a_215_47# 0.12fF
C6740 _390_/B _436_/a_68_297# 0.20fF
C6741 _459_/a_226_47# VPWR 0.08fF
C6742 _501_/a_109_47# _531_/A 0.23fF
C6743 _501_/a_397_297# _531_/C 0.12fF
C6744 _353_/X _419_/X 0.12fF
C6745 _442_/a_27_47# _478_/A 0.26fF
C6746 B[1] _383_/X 0.08fF
C6747 _390_/B output22/a_27_47# 0.19fF
C6748 _411_/A _481_/A 0.01fF
C6749 _375_/a_79_199# _376_/X 0.01fF
C6750 _328_/B _408_/B 0.13fF
C6751 VPWR _484_/a_215_47# 0.05fF
C6752 _406_/a_113_47# _406_/Y 0.08fF
C6753 _615_/a_78_199# _615_/a_215_47# 0.26fF
C6754 _448_/B _324_/a_62_47# 0.46fF
C6755 _557_/A _531_/C 0.27fF
C6756 _633_/Y _411_/A 0.60fF
C6757 _426_/A _432_/B 1.37fF
C6758 VPWR _531_/A 2.21fF
C6759 _516_/A _447_/B 1.32fF
C6760 _544_/A _542_/B 0.13fF
C6761 _567_/B _460_/a_489_413# 0.02fF
C6762 _549_/X _552_/a_489_413# 0.01fF
C6763 _562_/a_292_297# _627_/B 0.02fF
C6764 _386_/a_664_47# _480_/A 0.01fF
C6765 _613_/a_323_297# VPWR 0.02fF
C6766 input3/a_381_47# VPWR 0.33fF
C6767 _455_/X _359_/B 0.01fF
C6768 _385_/a_664_47# _385_/a_841_47# 0.29fF
C6769 _385_/a_62_47# _393_/A 0.55fF
C6770 input12/a_381_47# _442_/D 0.61fF
C6771 VPWR _469_/X 4.58fF
C6772 _455_/a_448_47# _418_/X 0.17fF
C6773 _551_/a_226_47# VPWR 0.09fF
C6774 _528_/a_384_47# _527_/A 0.09fF
C6775 _528_/a_81_21# _531_/B 0.24fF
C6776 _346_/a_161_47# _346_/A 0.58fF
C6777 _614_/a_489_413# _591_/A 0.02fF
C6778 _516_/A _376_/a_68_297# 0.00fF
C6779 _579_/a_59_75# _579_/X 0.30fF
C6780 _611_/X _621_/a_78_199# 0.33fF
C6781 _541_/a_292_297# _340_/A 0.01fF
C6782 _381_/C _485_/a_27_47# 0.28fF
C6783 _342_/X _417_/A 0.89fF
C6784 _455_/X _456_/a_76_199# 0.21fF
C6785 _546_/X _574_/a_81_21# 0.34fF
C6786 _471_/A _472_/B 0.21fF
C6787 _502_/a_292_297# VPWR 0.02fF
C6788 _338_/X _344_/a_215_47# 0.10fF
C6789 _391_/B _442_/B 0.28fF
C6790 _563_/a_109_297# _542_/D 0.01fF
C6791 _504_/a_227_47# _627_/A 0.11fF
C6792 _516_/A _386_/a_381_47# 0.12fF
C6793 _512_/a_78_199# VPWR 0.57fF
C6794 A[6] _547_/a_79_199# 0.04fF
C6795 _392_/A _406_/A 0.01fF
C6796 _430_/A _363_/A 0.04fF
C6797 _387_/a_493_297# _313_/A 0.08fF
C6798 _387_/a_78_199# _391_/A 0.23fF
C6799 VPWR M[3] 1.36fF
C6800 _501_/Y _531_/A 0.30fF
C6801 _576_/a_76_199# _574_/X 0.34fF
C6802 _576_/a_226_47# _575_/X 0.54fF
C6803 _386_/X _518_/a_256_47# 0.02fF
C6804 _330_/A B[5] 0.03fF
C6805 _443_/B _478_/A 0.04fF
C6806 _376_/X _419_/X 0.28fF
C6807 _603_/Y _553_/a_292_297# 0.08fF
C6808 VPWR _366_/a_76_199# 0.46fF
C6809 _410_/C _483_/X 0.36fF
C6810 _595_/X _598_/B 0.00fF
C6811 _491_/a_226_47# _489_/X 0.25fF
C6812 _427_/Y _427_/A 1.06fF
C6813 _407_/a_27_47# _406_/A 0.06fF
C6814 _407_/a_109_297# _406_/B 0.06fF
C6815 _440_/a_226_47# _440_/X 0.05fF
C6816 _520_/X _522_/a_489_413# 0.25fF
C6817 _464_/A VPWR 2.11fF
C6818 _586_/a_505_21# _503_/A 0.36fF
C6819 _510_/A _584_/A 0.06fF
C6820 _634_/Y _368_/a_68_297# 0.03fF
C6821 _349_/a_215_47# _350_/B 0.02fF
C6822 _543_/A _543_/Y 0.05fF
C6823 _570_/B _433_/Y 0.03fF
C6824 _381_/a_27_47# _381_/a_109_47# 0.03fF
C6825 _543_/B B[0] 0.53fF
C6826 _611_/X _627_/D 0.28fF
C6827 _419_/X _395_/X 0.13fF
C6828 _315_/a_161_47# VPWR 1.04fF
C6829 _404_/a_558_47# VPWR 0.36fF
C6830 _436_/A _351_/A 0.58fF
C6831 _613_/X _621_/X 0.39fF
C6832 _409_/a_78_199# _481_/A 0.37fF
C6833 _584_/A _485_/D 0.69fF
C6834 _545_/Y _588_/A 0.54fF
C6835 _607_/a_78_199# _606_/A 0.34fF
C6836 _328_/A _314_/a_68_297# 0.22fF
C6837 _347_/a_27_47# VPWR 0.83fF
C6838 _375_/X _384_/a_226_297# 0.01fF
C6839 _431_/X _428_/X 0.22fF
C6840 _432_/X _430_/X 0.43fF
C6841 input9/a_27_47# B[0] 0.37fF
C6842 _567_/B _521_/a_78_199# 0.00fF
C6843 _566_/A _565_/a_80_21# 0.20fF
C6844 _596_/a_76_199# _601_/A 0.01fF
C6845 _544_/A _563_/D 0.52fF
C6846 VPWR _546_/X 6.64fF
C6847 _566_/A _545_/Y 0.33fF
C6848 A[6] _410_/C 0.17fF
C6849 _631_/B VPWR 8.63fF
C6850 _569_/Y _572_/A 0.03fF
C6851 _417_/a_303_47# _542_/A 0.06fF
C6852 _563_/a_205_297# _627_/C 0.02fF
C6853 _535_/Y _539_/X 0.32fF
C6854 _469_/A _547_/X 0.03fF
C6855 _626_/Y _540_/X 0.28fF
C6856 _567_/Y _538_/Y 0.15fF
C6857 _406_/Y _433_/Y 0.35fF
C6858 _464_/A _501_/Y 0.04fF
C6859 input5/a_381_47# A[4] 0.02fF
C6860 B[0] _538_/Y 0.18fF
C6861 output29/a_27_47# _627_/B 0.10fF
C6862 _469_/A _570_/a_68_297# 0.02fF
C6863 _442_/a_303_47# VPWR 0.00fF
C6864 _327_/a_493_297# _481_/A 0.08fF
C6865 M[1] _633_/Y 0.04fF
C6866 _469_/a_381_47# _469_/a_841_47# 0.03fF
C6867 _563_/D _391_/B 1.85fF
C6868 _386_/A _510_/A 0.14fF
C6869 VPWR _411_/X 0.83fF
C6870 _370_/a_68_297# _370_/A 0.41fF
C6871 _561_/A _452_/a_68_297# 0.20fF
C6872 _468_/a_78_199# _468_/a_292_297# 0.03fF
C6873 _440_/X _439_/X 0.01fF
C6874 A[6] _507_/a_109_297# 0.02fF
C6875 VPWR _324_/a_841_47# 0.32fF
C6876 _429_/a_226_47# _432_/B 0.05fF
C6877 _607_/X _624_/X 0.03fF
C6878 _479_/B _486_/X 0.16fF
C6879 _447_/a_68_297# _447_/a_150_297# 0.02fF
C6880 _626_/Y _610_/Y 0.10fF
C6881 _506_/A _508_/a_77_199# 0.16fF
C6882 _374_/a_215_47# VPWR 0.08fF
C6883 _314_/X _631_/B 0.06fF
C6884 _433_/Y _381_/B 0.41fF
C6885 B[7] _452_/a_68_297# 0.08fF
C6886 _523_/a_76_199# VPWR 0.45fF
C6887 _351_/A _350_/X 0.02fF
C6888 _627_/D _622_/a_183_297# 0.01fF
C6889 _543_/A _585_/B 0.48fF
C6890 _463_/a_226_47# _497_/a_68_297# 0.01fF
C6891 _487_/X _515_/A 0.13fF
C6892 _567_/B _585_/B 0.53fF
C6893 _513_/A _479_/B 0.63fF
C6894 _536_/Y _587_/A 0.59fF
C6895 _544_/A _518_/a_250_297# 0.00fF
C6896 _602_/Y _558_/a_77_199# 0.01fF
C6897 _616_/B _624_/a_489_47# 0.02fF
C6898 _386_/A _485_/D 1.48fF
C6899 _488_/a_226_47# VPWR 0.07fF
C6900 _562_/a_292_297# VPWR 0.01fF
C6901 _392_/Y _406_/A 0.05fF
C6902 _525_/a_76_199# _525_/X 0.22fF
C6903 _559_/a_227_47# _570_/a_68_297# 0.04fF
C6904 _488_/a_76_199# _469_/A 0.07fF
C6905 _584_/A A[6] 0.05fF
C6906 _542_/A _484_/a_78_199# 0.01fF
C6907 _476_/a_93_21# _633_/Y 0.02fF
C6908 input6/a_27_47# _361_/a_226_47# 0.01fF
C6909 _444_/A _442_/B 0.10fF
C6910 _627_/A _533_/a_77_199# 0.05fF
C6911 _627_/D _627_/a_27_297# 0.32fF
C6912 _444_/A _542_/B 0.27fF
C6913 _531_/C _531_/A 2.17fF
C6914 _482_/a_68_297# VPWR 0.31fF
C6915 _381_/B _540_/X 0.03fF
C6916 _442_/B B[5] 0.03fF
C6917 _386_/a_664_47# _515_/Y 0.08fF
C6918 _544_/A _547_/a_222_93# 0.05fF
C6919 _487_/X _535_/Y 0.08fF
C6920 B[0] _486_/X 1.65fF
C6921 _371_/B _363_/B 2.93fF
C6922 _627_/X _627_/D 0.09fF
C6923 _455_/a_544_297# VPWR 0.01fF
C6924 _583_/X _633_/Y 0.02fF
C6925 _513_/A B[0] 0.03fF
C6926 _524_/a_78_199# _523_/X 0.06fF
C6927 _390_/D _313_/A 0.01fF
C6928 _521_/a_215_47# _488_/X 0.07fF
C6929 _451_/a_27_47# _584_/A 0.15fF
C6930 _613_/a_77_199# _613_/a_323_297# 0.05fF
C6931 _351_/X _361_/X 3.03fF
C6932 _571_/a_250_297# _570_/A 0.01fF
C6933 _570_/X _595_/X 0.00fF
C6934 _432_/a_68_297# _432_/X 0.27fF
C6935 _487_/a_78_199# _449_/A 0.23fF
C6936 _342_/X _631_/B 0.22fF
C6937 _555_/a_27_413# _554_/B 0.14fF
C6938 _375_/X _384_/X 0.27fF
C6939 _430_/A _426_/A 0.24fF
C6940 _378_/a_558_47# _378_/a_664_47# 0.60fF
C6941 _378_/a_381_47# _378_/a_841_47# 0.03fF
C6942 _386_/X _437_/a_222_93# 0.09fF
C6943 _442_/B _394_/a_558_47# 0.32fF
C6944 _521_/X _483_/X 0.01fF
C6945 _576_/a_226_297# _530_/X 0.01fF
C6946 _520_/X _503_/A 0.11fF
C6947 _386_/X _510_/A 0.03fF
C6948 _570_/A _515_/A 0.32fF
C6949 _456_/X _490_/a_292_297# 0.08fF
C6950 _378_/a_381_47# _367_/C 0.04fF
C6951 _457_/a_226_47# _456_/X 0.52fF
C6952 VPWR _548_/a_76_199# 0.45fF
C6953 _558_/a_77_199# _558_/a_227_297# 0.13fF
C6954 _567_/B _558_/X 0.03fF
C6955 _590_/A _503_/A 0.26fF
C6956 _436_/A _519_/A 0.14fF
C6957 _542_/C _515_/A 0.17fF
C6958 input15/a_75_212# _401_/A 0.22fF
C6959 _483_/a_93_21# _483_/X 0.13fF
C6960 _573_/Y _548_/a_489_413# 0.00fF
C6961 _544_/A _518_/X 0.33fF
C6962 _417_/A _351_/a_27_53# 0.09fF
C6963 _564_/A _572_/A 0.02fF
C6964 _497_/a_68_297# _498_/A 0.27fF
C6965 M[0] VPWR 0.84fF
C6966 _487_/a_493_297# _542_/A 0.02fF
C6967 _386_/A A[6] 0.16fF
C6968 _349_/a_493_297# VPWR 0.01fF
C6969 _511_/X _522_/a_76_199# 0.04fF
C6970 _519_/A _542_/D 0.07fF
C6971 _535_/Y _570_/A 0.60fF
C6972 _386_/X _485_/D 0.35fF
C6973 A[3] _539_/X 0.45fF
C6974 _410_/a_27_47# _442_/a_27_47# 0.01fF
C6975 _475_/X _633_/Y 0.64fF
C6976 _423_/X _363_/A 0.08fF
C6977 _446_/X _471_/A 0.56fF
C6978 _464_/A _531_/C 0.02fF
C6979 _433_/Y _542_/A 0.05fF
C6980 _500_/a_78_199# _465_/X 0.33fF
C6981 B[0] _451_/A 0.01fF
C6982 _569_/Y _589_/a_556_47# 0.02fF
C6983 _382_/a_68_297# VPWR 0.29fF
C6984 _469_/a_558_47# _610_/A 0.14fF
C6985 _543_/B _572_/A 0.24fF
C6986 _381_/C _381_/a_27_47# 0.19fF
C6987 A[6] _521_/X 0.00fF
C6988 _613_/a_539_297# _433_/Y 0.03fF
C6989 _567_/B _572_/B 0.06fF
C6990 _575_/X _485_/D 0.13fF
C6991 _515_/A _535_/A 0.50fF
C6992 _423_/a_78_199# _397_/a_489_413# 0.03fF
C6993 _371_/a_68_297# _430_/a_68_297# 0.00fF
C6994 _452_/a_68_297# VPWR 0.29fF
C6995 _557_/Y _602_/A 0.01fF
C6996 _483_/a_93_21# _483_/a_256_47# 0.03fF
C6997 _564_/A _542_/D 0.13fF
C6998 _375_/X _329_/a_76_199# 0.06fF
C6999 _613_/a_539_297# _586_/S 0.02fF
C7000 _613_/a_227_47# _612_/Y 0.19fF
C7001 _627_/A _469_/X 0.28fF
C7002 input3/a_664_47# _390_/D 0.05fF
C7003 A[6] _483_/a_93_21# 0.08fF
C7004 input5/a_558_47# _390_/B 0.08fF
C7005 _454_/a_226_47# _454_/X 0.15fF
C7006 _494_/a_226_297# _492_/X 0.03fF
C7007 _386_/X _483_/X 0.02fF
C7008 _467_/Y _557_/Y 0.16fF
C7009 _567_/B _533_/X 0.78fF
C7010 _404_/a_62_47# _469_/X 0.01fF
C7011 _633_/Y _574_/a_299_297# 0.18fF
C7012 _379_/a_292_297# _448_/B 0.02fF
C7013 _360_/a_76_199# _360_/a_489_413# 0.12fF
C7014 _386_/X _631_/A 0.02fF
C7015 _474_/A _503_/a_62_47# 0.02fF
C7016 _386_/a_664_47# _386_/a_841_47# 0.29fF
C7017 _591_/Y _591_/A 1.18fF
C7018 _626_/Y _494_/X 0.14fF
C7019 _386_/A _443_/A 0.13fF
C7020 _485_/A _481_/A 0.33fF
C7021 M[2] _343_/a_556_47# 0.02fF
C7022 VPWR output29/a_27_47# 0.64fF
C7023 _458_/a_292_297# VPWR 0.01fF
C7024 _535_/Y _535_/A 0.69fF
C7025 _326_/A _409_/a_215_47# 0.10fF
C7026 _543_/B _542_/D 0.16fF
C7027 _403_/a_27_47# _472_/B 0.31fF
C7028 _573_/Y _594_/X 0.56fF
C7029 M[7] _558_/a_227_47# 0.02fF
C7030 _400_/a_209_297# _631_/B 0.13fF
C7031 _530_/a_76_199# _529_/a_27_47# 0.00fF
C7032 _452_/X _453_/a_93_21# 0.09fF
C7033 _558_/a_77_199# _558_/X 0.26fF
C7034 _475_/X _475_/a_150_297# 0.01fF
C7035 _542_/B _482_/X 0.03fF
C7036 _378_/a_62_47# _324_/a_62_47# 0.02fF
C7037 _476_/X _525_/a_76_199# 0.01fF
C7038 _338_/a_448_47# VPWR 0.05fF
C7039 _544_/A _520_/X 0.04fF
C7040 _361_/a_76_199# _363_/B 0.00fF
C7041 _542_/a_27_47# _542_/A 0.43fF
C7042 _386_/X _483_/a_256_47# 0.03fF
C7043 _487_/X A[3] 0.11fF
C7044 _600_/a_285_47# VPWR 0.01fF
C7045 _619_/a_27_47# _607_/a_78_199# 0.00fF
C7046 _410_/a_27_47# _443_/B 0.20fF
C7047 _411_/B _442_/a_27_47# 0.01fF
C7048 _337_/A _320_/a_161_47# 0.07fF
C7049 _347_/A _350_/C 0.28fF
C7050 B[3] _618_/Y 0.00fF
C7051 _587_/a_27_47# _624_/a_206_369# 0.00fF
C7052 _597_/a_292_297# _559_/X 0.02fF
C7053 _386_/X A[6] 0.08fF
C7054 _597_/a_78_199# _576_/X 0.29fF
C7055 _435_/a_27_47# _587_/A 0.24fF
C7056 _632_/a_78_199# _632_/a_292_297# 0.03fF
C7057 _470_/a_80_21# _470_/a_209_47# 0.04fF
C7058 _459_/X _457_/X 1.35fF
C7059 _588_/A _622_/C 0.43fF
C7060 _595_/a_227_297# _588_/A 0.04fF
C7061 _430_/a_68_297# _432_/X 0.00fF
C7062 _607_/X _612_/A 0.05fF
C7063 _519_/X _484_/a_78_199# 0.12fF
C7064 _381_/C _382_/B 0.04fF
C7065 _587_/A _539_/A 2.64fF
C7066 _533_/a_227_47# VPWR 0.12fF
C7067 VPWR _462_/a_76_199# 0.61fF
C7068 _602_/Y _553_/a_78_199# 0.06fF
C7069 _633_/Y _367_/a_27_297# 0.02fF
C7070 _393_/A _363_/B 0.06fF
C7071 _445_/X _446_/a_250_297# 0.04fF
C7072 _417_/D _367_/C 1.49fF
C7073 _412_/a_489_413# _419_/X 0.13fF
C7074 _465_/a_27_297# _427_/Y 0.25fF
C7075 _568_/a_539_297# _566_/Y 0.03fF
C7076 _627_/C _541_/a_215_47# 0.01fF
C7077 _378_/A _542_/A 0.31fF
C7078 _478_/A _507_/Y 0.68fF
C7079 _347_/a_27_47# _563_/A 0.43fF
C7080 B[0] _627_/B 0.63fF
C7081 _557_/Y _606_/A 0.18fF
C7082 _603_/a_27_47# _555_/a_215_297# 0.04fF
C7083 _454_/X _453_/X 0.27fF
C7084 _602_/A _606_/A 0.19fF
C7085 _563_/A _631_/B 0.04fF
C7086 _332_/X _367_/C 0.20fF
C7087 _569_/Y _570_/B 0.19fF
C7088 _360_/a_489_413# _353_/X 0.07fF
C7089 _347_/A _442_/A 0.34fF
C7090 _493_/a_78_199# _460_/a_76_199# 0.04fF
C7091 _607_/X _625_/Y 0.03fF
C7092 B[7] _599_/Y 0.22fF
C7093 _404_/a_62_47# _404_/a_558_47# 0.03fF
C7094 _627_/A _546_/X 0.03fF
C7095 _461_/a_78_199# _390_/B 0.16fF
C7096 _469_/A _633_/Y 0.03fF
C7097 _607_/X _601_/Y 0.02fF
C7098 _567_/B _468_/a_215_47# 0.16fF
C7099 _382_/X _383_/a_226_47# 0.61fF
C7100 _366_/a_76_199# _368_/A 0.24fF
C7101 _534_/a_209_47# _485_/D 0.03fF
C7102 _494_/X _527_/A 0.01fF
C7103 _397_/X B[5] 0.03fF
C7104 _391_/A _419_/X 0.03fF
C7105 B[0] _561_/A 0.14fF
C7106 _485_/A _520_/a_556_47# 0.02fF
C7107 _467_/Y _427_/A 0.00fF
C7108 _424_/X _423_/X 0.72fF
C7109 A[3] _570_/A 0.03fF
C7110 _492_/a_489_413# _504_/X 0.11fF
C7111 _492_/a_76_199# _524_/X 0.01fF
C7112 _330_/A _384_/a_76_199# 0.01fF
C7113 _330_/A _351_/X 0.08fF
C7114 _550_/a_292_297# _522_/X 0.08fF
C7115 _548_/X _546_/X 0.09fF
C7116 B[0] B[7] 0.03fF
C7117 _411_/B _443_/B 0.76fF
C7118 _409_/a_78_199# _409_/a_292_297# 0.03fF
C7119 _376_/X _631_/A 0.00fF
C7120 _575_/X _598_/B 0.07fF
C7121 _630_/a_76_199# _630_/a_226_297# 0.01fF
C7122 _630_/a_226_47# _630_/a_489_413# 0.02fF
C7123 _617_/a_113_297# _618_/A 0.22fF
C7124 output25/a_27_47# _374_/a_215_47# 0.02fF
C7125 _468_/a_215_47# _468_/a_78_199# 0.26fF
C7126 _426_/B _426_/a_68_297# 0.30fF
C7127 _568_/a_77_199# _587_/A 0.02fF
C7128 _513_/A _542_/D 0.42fF
C7129 _509_/Y _511_/a_346_47# 0.04fF
C7130 _563_/D _482_/X 0.02fF
C7131 M[12] input12/a_381_47# 0.17fF
C7132 _623_/X _564_/a_219_297# 0.00fF
C7133 _547_/X _570_/a_68_297# 0.01fF
C7134 B[1] _481_/A 0.06fF
C7135 _448_/B _447_/B 1.03fF
C7136 _490_/X _489_/X 2.38fF
C7137 _591_/Y _590_/A 0.14fF
C7138 _554_/A _555_/a_215_297# 0.38fF
C7139 _534_/a_80_21# _386_/a_381_47# 0.03fF
C7140 _629_/A _371_/B 0.18fF
C7141 _633_/Y _489_/a_76_199# 0.08fF
C7142 _580_/A VPWR 1.92fF
C7143 _485_/a_27_47# _485_/D 0.21fF
C7144 _441_/a_215_47# _340_/A 0.05fF
C7145 _395_/X _631_/A 0.01fF
C7146 _500_/a_215_47# _467_/a_109_47# 0.00fF
C7147 _569_/Y _381_/B 0.21fF
C7148 _519_/a_111_297# _381_/C 0.03fF
C7149 _410_/a_109_47# _631_/Y 0.04fF
C7150 _454_/X _542_/D 0.07fF
C7151 _584_/A _590_/B 0.03fF
C7152 _382_/B _419_/X 0.63fF
C7153 _390_/D _472_/B 0.32fF
C7154 _355_/a_161_47# _322_/a_27_47# 0.04fF
C7155 _633_/A _475_/A 0.09fF
C7156 _533_/a_77_199# _533_/a_323_297# 0.05fF
C7157 _417_/D _380_/A 0.24fF
C7158 A[5] _330_/A 0.19fF
C7159 _396_/X _383_/X 0.11fF
C7160 _536_/Y _433_/Y 0.47fF
C7161 _433_/a_109_47# _433_/a_397_297# 0.05fF
C7162 _444_/Y _446_/X 0.02fF
C7163 _410_/B _443_/A 0.08fF
C7164 _390_/D _445_/a_68_297# 0.20fF
C7165 _609_/a_80_21# _609_/a_209_47# 0.04fF
C7166 _542_/B _487_/X 0.03fF
C7167 B[7] _454_/a_226_47# 0.07fF
C7168 _549_/a_76_199# _574_/X 0.01fF
C7169 _360_/X _445_/A 0.03fF
C7170 _408_/B _328_/A 1.93fF
C7171 _633_/A _633_/a_74_47# 0.47fF
C7172 _618_/A _601_/A 0.39fF
C7173 _616_/B _624_/X 0.03fF
C7174 _421_/a_76_199# _421_/a_226_47# 0.49fF
C7175 _615_/a_215_47# VPWR 0.17fF
C7176 _573_/A _590_/A 0.01fF
C7177 _513_/A _478_/A 0.07fF
C7178 _456_/X _454_/X 0.96fF
C7179 _587_/A _588_/A 1.23fF
C7180 _457_/X _504_/X 0.09fF
C7181 _451_/A _542_/D 0.82fF
C7182 _383_/X _481_/A 1.17fF
C7183 _479_/B VPWR 1.52fF
C7184 _324_/a_558_47# _324_/a_841_47# 0.07fF
C7185 _612_/A _588_/A 0.10fF
C7186 _322_/A _441_/a_78_199# 0.01fF
C7187 _623_/X _442_/D 0.11fF
C7188 _583_/X _625_/a_27_297# 0.14fF
C7189 _474_/A _510_/X 0.16fF
C7190 _445_/A _409_/a_215_47# 0.12fF
C7191 _550_/X _522_/X 0.01fF
C7192 _356_/a_215_47# _481_/A 0.10fF
C7193 _633_/Y _383_/X 0.07fF
C7194 _566_/A _587_/A 0.03fF
C7195 _598_/a_68_297# VPWR 0.28fF
C7196 _471_/Y _503_/A 0.41fF
C7197 _452_/A _449_/A 0.01fF
C7198 _454_/X _346_/A 0.20fF
C7199 _504_/a_227_47# _468_/a_78_199# 0.07fF
C7200 _341_/a_27_47# _436_/A 0.50fF
C7201 VPWR _599_/Y 1.50fF
C7202 _578_/a_215_47# _550_/X 0.11fF
C7203 input5/a_62_47# VPWR 0.51fF
C7204 _454_/X _478_/A 0.07fF
C7205 _583_/X _616_/Y 2.09fF
C7206 _530_/X _486_/a_68_297# 0.15fF
C7207 _502_/a_493_297# _494_/X 0.04fF
C7208 _502_/a_215_47# _468_/X 0.03fF
C7209 _541_/a_78_199# _514_/A 0.01fF
C7210 _386_/X _446_/a_250_297# 0.03fF
C7211 _583_/X _563_/B 0.01fF
C7212 _567_/B _557_/A 0.40fF
C7213 _544_/a_558_47# _588_/A 0.11fF
C7214 _362_/a_76_199# _363_/B 0.22fF
C7215 _623_/X _588_/Y 0.31fF
C7216 _625_/Y _588_/A 0.34fF
C7217 _485_/a_27_47# A[6] 0.10fF
C7218 _567_/Y VPWR 1.60fF
C7219 _620_/X _625_/a_27_47# 0.01fF
C7220 _447_/X output32/a_27_47# 0.01fF
C7221 _532_/a_206_369# _528_/a_299_297# 0.00fF
C7222 _561_/A _453_/X 0.00fF
C7223 _519_/X _378_/A 0.09fF
C7224 _424_/a_76_199# _424_/a_489_413# 0.12fF
C7225 B[0] VPWR 2.55fF
C7226 _351_/X _442_/B 0.46fF
C7227 _375_/X _328_/A 0.69fF
C7228 _444_/Y _442_/D 0.24fF
C7229 _395_/X _391_/a_68_297# 0.03fF
C7230 _351_/a_219_297# _363_/B 0.01fF
C7231 _542_/B _570_/A 0.03fF
C7232 _548_/a_76_199# _548_/X 0.22fF
C7233 _626_/a_109_297# _623_/X 0.01fF
C7234 VPWR _521_/a_292_297# 0.01fF
C7235 _626_/a_109_47# _625_/Y 0.54fF
C7236 _620_/X _616_/A 0.54fF
C7237 _572_/A _627_/B 0.36fF
C7238 B[7] _453_/X 0.68fF
C7239 _542_/C _442_/B 0.73fF
C7240 _604_/a_80_21# _558_/a_227_47# 0.06fF
C7241 M[2] _634_/a_384_47# 0.01fF
C7242 _491_/X _492_/a_76_199# 0.22fF
C7243 _476_/X _492_/a_226_47# 0.27fF
C7244 _628_/a_28_47# _628_/a_300_47# 0.50fF
C7245 _436_/A _395_/a_150_297# 0.01fF
C7246 _542_/B _542_/C 4.40fF
C7247 _469_/A _521_/a_78_199# 0.09fF
C7248 _408_/X VPWR 1.52fF
C7249 VPWR _468_/a_493_297# 0.01fF
C7250 _622_/a_29_53# _627_/B 0.61fF
C7251 VPWR _320_/a_161_47# 0.97fF
C7252 output18/a_27_47# M[10] 0.46fF
C7253 _343_/a_489_413# _338_/X 0.25fF
C7254 _584_/A _394_/a_664_47# 0.05fF
C7255 _336_/a_78_199# _367_/C 0.33fF
C7256 _536_/Y _537_/a_539_297# 0.02fF
C7257 _566_/Y _503_/A 0.14fF
C7258 _461_/X _460_/X 1.40fF
C7259 _506_/A _483_/X 0.31fF
C7260 _396_/a_93_21# _631_/B 0.11fF
C7261 _423_/a_215_47# _631_/A 0.16fF
C7262 _379_/a_215_47# _417_/A 0.35fF
C7263 _608_/a_78_199# _627_/B 0.53fF
C7264 B[7] _616_/A 0.11fF
C7265 _538_/Y _570_/B 0.00fF
C7266 _476_/a_93_21# _476_/a_250_297# 0.50fF
C7267 _630_/a_226_47# _629_/a_68_297# 0.00fF
C7268 _419_/X _421_/a_76_199# 0.29fF
C7269 _487_/X _563_/D 0.03fF
C7270 _455_/X _347_/A 0.55fF
C7271 _492_/X VPWR 1.58fF
C7272 _605_/a_80_21# _557_/Y 0.03fF
C7273 _338_/a_79_199# _366_/a_226_47# 0.01fF
C7274 _629_/X _432_/B 1.27fF
C7275 _582_/a_27_47# VPWR 0.03fF
C7276 _552_/a_76_199# _552_/a_226_47# 0.49fF
C7277 _542_/D _627_/B 0.41fF
C7278 _583_/a_556_47# VPWR 0.01fF
C7279 _365_/a_299_297# _630_/X 0.00fF
C7280 _454_/a_226_47# VPWR 0.23fF
C7281 _628_/a_300_47# _622_/X 0.19fF
C7282 _523_/a_76_199# _523_/X 0.32fF
C7283 VPWR _344_/a_78_199# 0.81fF
C7284 _410_/B _446_/a_250_297# 0.07fF
C7285 _448_/a_150_297# _542_/D 0.01fF
C7286 _455_/a_448_47# _419_/a_226_47# 0.03fF
C7287 _578_/a_215_47# _530_/X 0.02fF
C7288 _620_/a_226_47# _620_/X 0.05fF
C7289 _620_/a_489_413# _618_/Y 0.07fF
C7290 _381_/B _507_/Y 0.11fF
C7291 _629_/A _393_/A 0.02fF
C7292 _386_/A _388_/a_27_47# 0.12fF
C7293 VPWR _558_/a_323_297# 0.02fF
C7294 _557_/A _558_/a_77_199# 0.30fF
C7295 _390_/a_27_47# _391_/B 0.20fF
C7296 _487_/X _477_/a_292_297# 0.02fF
C7297 _419_/X _442_/B 0.75fF
C7298 _352_/X VPWR 2.33fF
C7299 _553_/a_78_199# _553_/a_292_297# 0.03fF
C7300 A[3] _621_/X 0.03fF
C7301 _469_/A _585_/B 0.19fF
C7302 _506_/A A[6] 1.05fF
C7303 _436_/X _390_/B 0.31fF
C7304 _352_/X _361_/a_226_297# 0.02fF
C7305 _485_/D _515_/A 0.72fF
C7306 _530_/X _486_/B 0.10fF
C7307 _448_/B _418_/X 0.04fF
C7308 _561_/A _542_/D 2.21fF
C7309 _510_/A _385_/a_664_47# 0.12fF
C7310 _613_/X _590_/B 0.02fF
C7311 _627_/A _533_/a_227_47# 0.31fF
C7312 _485_/A _563_/B 0.02fF
C7313 _567_/B _527_/Y 0.04fF
C7314 _338_/a_222_93# _631_/B 0.08fF
C7315 _572_/B _574_/a_299_297# 0.07fF
C7316 _572_/A _574_/a_81_21# 0.20fF
C7317 _337_/a_68_297# _337_/B 0.30fF
C7318 B[7] _542_/D 0.16fF
C7319 _418_/B M[9] 0.05fF
C7320 _350_/C _410_/C 0.15fF
C7321 _471_/Y _504_/X 0.01fF
C7322 _433_/Y _539_/A 0.31fF
C7323 _313_/A _313_/a_27_47# 0.40fF
C7324 _485_/D _535_/Y 0.37fF
C7325 _417_/D _452_/A 0.70fF
C7326 _563_/D _570_/A 0.05fF
C7327 _538_/Y _381_/B 0.13fF
C7328 _448_/A _453_/a_250_297# 0.06fF
C7329 _440_/X _460_/X 0.43fF
C7330 _360_/X _371_/B 0.03fF
C7331 _577_/a_76_199# _390_/D 0.07fF
C7332 _476_/a_250_297# _475_/X 0.29fF
C7333 _346_/a_161_47# _340_/a_27_47# 0.03fF
C7334 _365_/a_299_297# _363_/B 0.19fF
C7335 _347_/A _477_/a_215_47# 0.18fF
C7336 _448_/a_68_297# _448_/B 0.30fF
C7337 _493_/a_292_297# _458_/X 0.06fF
C7338 _544_/A _566_/Y 0.04fF
C7339 _611_/X _623_/X 0.88fF
C7340 _386_/a_381_47# _514_/B 0.01fF
C7341 _338_/a_448_47# _368_/A 0.07fF
C7342 _338_/a_79_199# _337_/X 0.27fF
C7343 _519_/A _542_/A 0.70fF
C7344 _417_/A _363_/A 0.65fF
C7345 _627_/C _622_/X 0.01fF
C7346 _474_/Y _503_/A 0.23fF
C7347 _615_/a_78_199# _593_/A 0.12fF
C7348 _453_/X VPWR 1.15fF
C7349 _587_/A _616_/B 0.08fF
C7350 _417_/A _420_/X 2.93fF
C7351 _334_/a_303_47# VPWR 0.01fF
C7352 _612_/A _616_/B 0.38fF
C7353 _369_/a_76_199# _369_/a_226_47# 0.49fF
C7354 _360_/X _361_/a_489_413# 0.26fF
C7355 VPWR _625_/a_27_47# 0.05fF
C7356 _605_/a_80_21# _606_/A 0.31fF
C7357 _539_/A _540_/X 0.01fF
C7358 _604_/X M[7] 0.50fF
C7359 _474_/A _473_/a_77_199# 0.22fF
C7360 _620_/X _619_/Y 0.01fF
C7361 output17/a_27_47# _552_/a_226_47# 0.02fF
C7362 _336_/a_215_47# _332_/X 0.16fF
C7363 _442_/A _410_/C 0.21fF
C7364 _469_/a_381_47# _545_/Y 0.12fF
C7365 _474_/A _390_/B 0.06fF
C7366 _422_/X VPWR 3.00fF
C7367 _633_/Y _547_/X 0.11fF
C7368 _603_/Y M[0] 0.00fF
C7369 _523_/a_489_413# _631_/Y 0.11fF
C7370 _385_/a_558_47# _475_/A 0.08fF
C7371 _510_/A _391_/A 0.20fF
C7372 _634_/a_27_413# _634_/a_300_297# 0.04fF
C7373 _625_/Y _625_/a_277_47# 0.24fF
C7374 _417_/D _540_/a_250_297# 0.09fF
C7375 _390_/D _446_/X 0.52fF
C7376 _580_/B _581_/B 0.01fF
C7377 VPWR _616_/A 5.09fF
C7378 VPWR _409_/a_493_297# 0.01fF
C7379 _342_/X _344_/a_78_199# 0.27fF
C7380 _599_/A _625_/a_27_297# 0.00fF
C7381 _619_/a_27_47# _606_/A 0.00fF
C7382 _381_/C _547_/a_222_93# 0.13fF
C7383 _579_/X _555_/a_215_297# 0.01fF
C7384 _567_/B _459_/a_226_47# 0.13fF
C7385 _418_/a_68_297# VPWR 0.29fF
C7386 _631_/Y _472_/B 0.03fF
C7387 _610_/A _624_/a_76_199# 0.07fF
C7388 _625_/Y _616_/B 0.94fF
C7389 _607_/X _610_/Y 0.07fF
C7390 _381_/B _486_/X 0.26fF
C7391 _518_/a_250_297# _570_/A 0.14fF
C7392 _336_/a_493_297# _442_/B 0.02fF
C7393 _398_/a_489_413# _399_/a_78_199# 0.02fF
C7394 _412_/X _420_/X 0.06fF
C7395 _429_/a_76_199# _350_/X 0.35fF
C7396 _584_/A _350_/C 1.12fF
C7397 _542_/A _507_/Y 0.11fF
C7398 _382_/A _382_/B 0.19fF
C7399 _475_/X _468_/a_215_47# 0.01fF
C7400 _572_/A VPWR 3.26fF
C7401 _396_/a_93_21# _396_/a_256_47# 0.03fF
C7402 _599_/A _616_/Y 0.03fF
C7403 _543_/B _542_/A 0.49fF
C7404 _601_/Y _616_/B 0.01fF
C7405 _442_/A _507_/a_109_297# 0.02fF
C7406 _487_/X _518_/X 0.03fF
C7407 _563_/D _419_/X 0.14fF
C7408 _568_/a_77_199# _433_/Y 0.06fF
C7409 _513_/A _381_/B 0.49fF
C7410 _580_/a_68_297# _580_/a_150_297# 0.02fF
C7411 VPWR _622_/a_29_53# 0.37fF
C7412 _520_/X _539_/X 0.49fF
C7413 _410_/B _506_/Y 0.03fF
C7414 _567_/B _469_/X 0.17fF
C7415 _590_/B _590_/a_68_297# 0.64fF
C7416 _338_/X _442_/B 0.03fF
C7417 _436_/A VPWR 5.70fF
C7418 _551_/X VPWR 1.21fF
C7419 _351_/A _363_/B 0.03fF
C7420 _608_/a_78_199# VPWR 0.62fF
C7421 _480_/Y _505_/a_80_21# 0.31fF
C7422 M[13] _626_/a_397_297# 0.01fF
C7423 _620_/a_226_47# VPWR 0.09fF
C7424 _476_/a_346_47# _587_/A 0.05fF
C7425 _375_/X _397_/a_226_47# 0.00fF
C7426 _381_/C _518_/X 0.16fF
C7427 _454_/X _381_/B 0.14fF
C7428 _584_/A _442_/A 0.03fF
C7429 _359_/X _383_/X 0.10fF
C7430 _474_/A _471_/A 0.08fF
C7431 _474_/Y _471_/Y 0.47fF
C7432 VPWR _542_/D 8.93fF
C7433 _631_/Y _554_/A 0.03fF
C7434 _359_/a_68_297# _359_/A 0.35fF
C7435 _482_/X _483_/a_250_297# 0.04fF
C7436 _448_/a_68_297# _453_/a_93_21# 0.01fF
C7437 B[2] _597_/a_215_47# 0.08fF
C7438 _390_/D _442_/D 0.12fF
C7439 _380_/A _410_/C 0.17fF
C7440 _627_/X _623_/X 0.23fF
C7441 _511_/a_346_47# _469_/X 0.10fF
C7442 _505_/a_209_47# _481_/A 0.07fF
C7443 _381_/a_27_47# A[6] 0.06fF
C7444 _461_/a_78_199# _406_/B 0.01fF
C7445 _349_/a_215_47# _351_/A 0.14fF
C7446 _465_/a_27_297# _427_/A 0.37fF
C7447 _417_/D _479_/a_68_297# 0.15fF
C7448 _504_/a_77_199# _436_/X 0.00fF
C7449 _331_/a_27_47# _384_/a_76_199# 0.02fF
C7450 _588_/A _433_/Y 0.17fF
C7451 _518_/X _570_/A 0.05fF
C7452 _360_/X _361_/a_76_199# 0.24fF
C7453 _623_/a_76_199# _623_/a_489_413# 0.12fF
C7454 _456_/X VPWR 2.35fF
C7455 VPWR _553_/a_493_297# 0.01fF
C7456 A[3] _485_/D 0.03fF
C7457 _417_/A _329_/X 0.37fF
C7458 _396_/a_250_297# _396_/X 0.03fF
C7459 M[11] VPWR 0.53fF
C7460 _429_/a_226_47# _429_/a_489_413# 0.02fF
C7461 _429_/a_76_199# _429_/a_226_297# 0.01fF
C7462 _612_/Y _588_/Y 0.71fF
C7463 _347_/A _541_/a_78_199# 0.15fF
C7464 _586_/S _588_/A 0.26fF
C7465 VPWR _350_/X 3.30fF
C7466 _566_/A _433_/Y 0.02fF
C7467 _475_/X _504_/a_227_47# 0.05fF
C7468 _487_/X _520_/X 1.85fF
C7469 A[5] _397_/X 0.06fF
C7470 _567_/Y _627_/A 0.03fF
C7471 _386_/X _406_/A 0.36fF
C7472 _423_/X _383_/X 0.01fF
C7473 _422_/a_226_47# _422_/a_489_413# 0.02fF
C7474 _422_/a_76_199# _422_/a_226_297# 0.01fF
C7475 _587_/A _530_/X 0.03fF
C7476 VPWR _346_/A 1.69fF
C7477 _469_/A _595_/a_227_47# 0.05fF
C7478 B[0] _627_/A 0.05fF
C7479 _610_/A _584_/A 0.55fF
C7480 _404_/a_558_47# _543_/A 0.14fF
C7481 _410_/C _316_/a_381_47# 0.69fF
C7482 _500_/a_493_297# _464_/A 0.13fF
C7483 VPWR _478_/A 5.03fF
C7484 _542_/A _486_/X 0.30fF
C7485 _588_/A _540_/X 0.24fF
C7486 VPWR _369_/a_489_413# 0.33fF
C7487 _386_/A _442_/A 0.03fF
C7488 A[3] _483_/X 0.73fF
C7489 input13/a_27_47# B[4] 0.38fF
C7490 _619_/Y VPWR 1.03fF
C7491 _477_/a_78_199# _477_/a_215_47# 0.26fF
C7492 _444_/A _446_/a_93_21# 0.02fF
C7493 _543_/Y _547_/X 0.27fF
C7494 _515_/Y _547_/X 0.27fF
C7495 _519_/X _520_/a_489_413# 0.14fF
C7496 _343_/a_76_199# _343_/X 0.29fF
C7497 _567_/B _546_/X 1.40fF
C7498 _525_/a_76_199# _525_/a_226_297# 0.01fF
C7499 _525_/a_226_47# _525_/a_489_413# 0.02fF
C7500 _519_/X _519_/A 0.15fF
C7501 _513_/A _542_/A 3.06fF
C7502 _626_/Y _620_/X 0.10fF
C7503 _330_/A _631_/A 1.11fF
C7504 _524_/a_215_47# _524_/X 0.03fF
C7505 _380_/A _584_/A 1.18fF
C7506 _448_/A _449_/A 0.20fF
C7507 _391_/A _391_/a_68_297# 0.30fF
C7508 _606_/Y _619_/Y 0.40fF
C7509 _433_/a_109_47# VPWR 0.25fF
C7510 _373_/a_199_47# _371_/A 0.15fF
C7511 _373_/a_113_297# _371_/B 0.09fF
C7512 _338_/a_222_93# _338_/a_448_47# 0.03fF
C7513 _422_/a_76_199# _421_/X 0.22fF
C7514 _426_/B _432_/X 0.01fF
C7515 _614_/a_76_199# _612_/Y 0.07fF
C7516 _474_/A _504_/a_77_199# 0.00fF
C7517 _576_/a_76_199# _576_/a_226_47# 0.49fF
C7518 _610_/Y _588_/A 0.41fF
C7519 _417_/D _538_/A 0.08fF
C7520 _423_/X _407_/Y 0.12fF
C7521 _626_/Y B[7] 0.73fF
C7522 _390_/B _431_/X 0.43fF
C7523 _454_/X _542_/A 1.76fF
C7524 _420_/X _631_/B 2.66fF
C7525 _604_/a_209_297# _557_/B 0.09fF
C7526 _591_/Y _573_/A 0.37fF
C7527 _569_/A _595_/X 0.21fF
C7528 _378_/A _340_/A 0.06fF
C7529 _340_/A _346_/a_161_47# 0.16fF
C7530 _408_/B _313_/a_27_47# 0.32fF
C7531 _632_/a_78_199# _631_/A 0.01fF
C7532 _336_/a_78_199# _336_/a_215_47# 0.26fF
C7533 _602_/A _556_/A 0.36fF
C7534 _520_/X _570_/A 0.90fF
C7535 _442_/D _389_/a_27_47# 0.38fF
C7536 _557_/Y _556_/A 0.71fF
C7537 _626_/a_109_47# _610_/Y 0.05fF
C7538 A[6] A[3] 0.67fF
C7539 _318_/a_27_47# _381_/C 0.37fF
C7540 _542_/C _520_/X 0.03fF
C7541 _455_/X _410_/C 0.05fF
C7542 _570_/X _571_/a_250_297# 0.28fF
C7543 _440_/X _493_/X 0.01fF
C7544 _563_/B _484_/a_493_297# 0.12fF
C7545 _518_/a_93_21# _518_/a_346_47# 0.05fF
C7546 _358_/a_109_47# _442_/A 0.01fF
C7547 _499_/a_81_21# _467_/Y 0.12fF
C7548 _404_/a_381_47# _585_/B 0.02fF
C7549 _479_/A _505_/a_80_21# 0.01fF
C7550 _442_/D _316_/a_558_47# 0.23fF
C7551 _510_/A _442_/B 0.24fF
C7552 _479_/B _505_/a_209_297# 0.03fF
C7553 _445_/A _313_/A 0.55fF
C7554 _430_/A _432_/B 0.14fF
C7555 _489_/a_226_47# _489_/a_489_413# 0.02fF
C7556 _423_/a_78_199# VPWR 0.63fF
C7557 B[2] _583_/X 0.08fF
C7558 _313_/A _395_/a_68_297# 0.00fF
C7559 _629_/A _365_/a_299_297# 0.05fF
C7560 _607_/a_78_199# _607_/a_292_297# 0.03fF
C7561 _480_/A _481_/A 0.95fF
C7562 _493_/a_78_199# VPWR 0.59fF
C7563 _322_/A _381_/C 0.10fF
C7564 _386_/X _442_/A 0.03fF
C7565 _585_/B _547_/X 0.22fF
C7566 _447_/a_68_297# _418_/B 0.00fF
C7567 _423_/a_493_297# _384_/X 0.02fF
C7568 _367_/a_27_297# _367_/a_109_297# 0.02fF
C7569 _417_/D _488_/X 0.35fF
C7570 _503_/A _539_/X 0.95fF
C7571 _556_/Y _604_/a_209_297# 0.24fF
C7572 _604_/X _604_/a_80_21# 0.22fF
C7573 _384_/a_489_413# _384_/a_76_199# 0.12fF
C7574 _520_/X _535_/A 0.04fF
C7575 _328_/X _631_/B 0.16fF
C7576 output31/a_27_47# VPWR 0.64fF
C7577 _533_/a_227_297# _539_/A 0.04fF
C7578 _347_/A _475_/A 0.10fF
C7579 _342_/X _369_/a_489_413# 0.07fF
C7580 _411_/A _411_/X 0.03fF
C7581 _613_/a_77_199# _622_/a_29_53# 0.03fF
C7582 _487_/a_215_47# _453_/X 0.20fF
C7583 _542_/B _485_/D 0.03fF
C7584 _611_/X _612_/Y 0.48fF
C7585 _506_/A _506_/Y 0.47fF
C7586 _469_/a_381_47# _622_/C 0.05fF
C7587 _570_/X _535_/Y 0.01fF
C7588 _588_/a_109_297# _627_/D 0.02fF
C7589 _390_/D _576_/X 0.36fF
C7590 _528_/a_384_47# _530_/X 0.05fF
C7591 _593_/Y _601_/A 0.25fF
C7592 _547_/a_79_199# _547_/a_448_47# 0.13fF
C7593 _350_/X _399_/a_215_47# 0.03fF
C7594 _418_/A _378_/a_381_47# 0.18fF
C7595 _410_/B _350_/C 0.08fF
C7596 _417_/A output32/a_27_47# 0.02fF
C7597 _533_/X _551_/a_76_199# 0.07fF
C7598 _633_/Y _481_/A 0.59fF
C7599 _455_/X _584_/A 0.03fF
C7600 _536_/Y _538_/Y 0.02fF
C7601 output21/a_27_47# _620_/X 0.47fF
C7602 _559_/X _540_/X 1.19fF
C7603 _397_/X _398_/X 1.10fF
C7604 _440_/a_489_413# _436_/X 0.16fF
C7605 _518_/a_584_47# _517_/X 0.03fF
C7606 _442_/B _631_/A 0.29fF
C7607 _612_/Y _618_/A 0.60fF
C7608 _390_/D _618_/A 0.00fF
C7609 _503_/a_381_47# _446_/X 0.12fF
C7610 _476_/a_93_21# _469_/X 0.32fF
C7611 _570_/B VPWR 2.91fF
C7612 output31/a_27_47# _501_/Y 0.44fF
C7613 _626_/Y VPWR 4.12fF
C7614 _524_/a_493_297# _490_/X 0.08fF
C7615 _524_/a_215_47# _491_/X 0.20fF
C7616 _410_/B _442_/A 1.17fF
C7617 _360_/X _362_/a_76_199# 0.09fF
C7618 _487_/X _503_/A 0.18fF
C7619 _613_/X _610_/A 0.36fF
C7620 _586_/a_76_199# _586_/a_505_21# 0.02fF
C7621 _498_/Y _468_/X 0.01fF
C7622 _495_/a_489_413# _492_/X 0.02fF
C7623 _488_/a_489_413# _486_/X 0.07fF
C7624 _627_/A _572_/A 0.19fF
C7625 A[1] _558_/X 0.46fF
C7626 _520_/a_76_199# _547_/a_79_199# 0.01fF
C7627 _436_/A _563_/A 0.66fF
C7628 VPWR _467_/a_109_47# 0.23fF
C7629 _544_/A _378_/a_664_47# 0.05fF
C7630 _374_/a_215_47# _374_/X 0.01fF
C7631 _513_/A _519_/X 0.26fF
C7632 _431_/a_489_413# _428_/X 0.07fF
C7633 _540_/a_250_297# _410_/C 0.04fF
C7634 _404_/a_62_47# _572_/A 0.14fF
C7635 _542_/B A[6] 0.05fF
C7636 _563_/D _510_/A 0.05fF
C7637 _610_/Y _625_/a_277_47# 0.01fF
C7638 _383_/a_76_199# VPWR 0.51fF
C7639 _442_/D _631_/Y 0.32fF
C7640 _563_/A _542_/D 0.39fF
C7641 _503_/A _438_/X 0.68fF
C7642 _610_/A _609_/a_80_21# 0.20fF
C7643 _406_/Y VPWR 2.47fF
C7644 _608_/a_292_297# _586_/S 0.02fF
C7645 _390_/D _549_/X 0.22fF
C7646 _579_/X _631_/Y 0.01fF
C7647 _375_/X _376_/a_68_297# 0.00fF
C7648 _519_/A _328_/a_68_297# 0.00fF
C7649 _417_/A _485_/A 0.02fF
C7650 _608_/a_78_199# _627_/A 0.01fF
C7651 _572_/B _547_/X 0.11fF
C7652 _455_/X _386_/A 0.03fF
C7653 _554_/X _602_/A 0.50fF
C7654 _490_/a_78_199# _446_/X 0.33fF
C7655 _457_/a_76_199# _446_/X 0.19fF
C7656 _554_/X _557_/Y 0.32fF
C7657 _516_/A _379_/a_493_297# 0.08fF
C7658 _514_/a_68_297# _514_/B 0.33fF
C7659 _561_/A _542_/A 1.95fF
C7660 _360_/X _374_/a_78_199# 0.13fF
C7661 M[8] _467_/a_481_47# 0.01fF
C7662 _610_/Y _616_/B 0.12fF
C7663 _385_/a_62_47# VPWR 0.48fF
C7664 B[7] _593_/A 0.03fF
C7665 _563_/D _485_/D 0.05fF
C7666 _627_/A _542_/D 0.37fF
C7667 _420_/a_79_199# _452_/A 0.12fF
C7668 _626_/Y _501_/Y 0.05fF
C7669 _569_/A _584_/A 0.05fF
C7670 _516_/A _520_/a_489_413# 0.11fF
C7671 _516_/A _519_/A 0.49fF
C7672 _600_/a_27_297# _599_/Y 0.14fF
C7673 B[7] _542_/A 0.17fF
C7674 _386_/X _316_/a_381_47# 0.16fF
C7675 _347_/A _390_/B 0.03fF
C7676 _613_/a_539_297# B[7] 0.04fF
C7677 VPWR _381_/B 4.18fF
C7678 _343_/a_76_199# _370_/B 0.00fF
C7679 _475_/X _469_/X 0.13fF
C7680 _525_/a_489_413# _492_/a_489_413# 0.02fF
C7681 _563_/A _350_/X 0.17fF
C7682 _503_/A _570_/A 0.29fF
C7683 _443_/A _442_/B 0.00fF
C7684 _371_/A _431_/X 0.09fF
C7685 _436_/A _351_/a_27_53# 0.01fF
C7686 _629_/B _432_/X 0.65fF
C7687 _417_/D _418_/A 0.87fF
C7688 output28/a_27_47# VPWR 0.41fF
C7689 _394_/a_381_47# _394_/a_664_47# 0.09fF
C7690 _460_/X _462_/a_226_297# 0.03fF
C7691 _496_/a_215_47# _406_/Y 0.20fF
C7692 _520_/X _540_/a_93_21# 0.09fF
C7693 _593_/A _574_/a_81_21# 0.01fF
C7694 _360_/a_76_199# _455_/X 0.26fF
C7695 _527_/A VPWR 1.97fF
C7696 _416_/a_78_199# _367_/C 0.03fF
C7697 _524_/X _554_/B 0.01fF
C7698 _353_/X _375_/a_222_93# 0.03fF
C7699 _584_/A _627_/D 0.85fF
C7700 _570_/X A[3] 0.16fF
C7701 _469_/a_381_47# _587_/A 0.12fF
C7702 _576_/a_76_199# _485_/D 0.07fF
C7703 _410_/B _380_/A 0.23fF
C7704 _569_/Y _588_/A 0.56fF
C7705 _559_/a_77_199# _535_/Y 0.20fF
C7706 _544_/A _487_/X 0.20fF
C7707 _523_/a_226_297# _511_/X 0.02fF
C7708 _523_/a_489_413# _522_/X 0.14fF
C7709 _478_/a_27_47# _479_/B 0.18fF
C7710 _337_/A _337_/X 0.36fF
C7711 _590_/A _621_/X 0.22fF
C7712 _610_/A _590_/a_68_297# 0.14fF
C7713 _485_/A _484_/a_215_47# 0.01fF
C7714 output25/a_27_47# _369_/a_489_413# 0.01fF
C7715 _539_/A _507_/Y 1.02fF
C7716 _393_/A input14/a_27_47# 0.22fF
C7717 _627_/A _478_/A 1.01fF
C7718 _569_/Y _566_/A 0.56fF
C7719 _497_/A _467_/Y 2.02fF
C7720 _410_/a_27_47# VPWR 0.83fF
C7721 M[9] _367_/C 0.03fF
C7722 output24/a_27_47# _588_/Y 0.00fF
C7723 _479_/a_68_297# _410_/C 0.01fF
C7724 _610_/Y _592_/a_113_297# 0.00fF
C7725 output21/a_27_47# VPWR 0.64fF
C7726 _469_/a_62_47# VPWR 0.51fF
C7727 _433_/Y _530_/X 0.02fF
C7728 B[2] _599_/A 0.83fF
C7729 _454_/a_226_297# _628_/Y 0.01fF
C7730 _355_/A _442_/D 0.15fF
C7731 _404_/a_381_47# _608_/X 0.01fF
C7732 _633_/A _632_/a_215_47# 0.01fF
C7733 _455_/X _386_/X 0.03fF
C7734 _473_/a_227_297# _472_/B 0.02fF
C7735 _425_/a_226_297# _407_/Y 0.04fF
C7736 _544_/A _381_/C 0.03fF
C7737 _385_/a_558_47# _394_/a_841_47# 0.01fF
C7738 _328_/B _332_/X 0.41fF
C7739 _445_/A _408_/B 0.28fF
C7740 _563_/D A[6] 0.08fF
C7741 _351_/a_27_53# _350_/X 0.20fF
C7742 _542_/C _390_/a_27_47# 0.32fF
C7743 _633_/Y _521_/a_78_199# 0.15fF
C7744 _408_/B _395_/a_68_297# 0.06fF
C7745 _546_/a_76_199# _546_/a_489_413# 0.12fF
C7746 B[0] _540_/a_584_47# 0.01fF
C7747 _538_/Y _539_/A 0.09fF
C7748 _530_/X _540_/X 0.03fF
C7749 _489_/a_226_47# _483_/X 0.16fF
C7750 _527_/B _532_/a_205_47# 0.08fF
C7751 _501_/a_109_297# _531_/A 0.01fF
C7752 _459_/a_489_413# VPWR 0.39fF
C7753 _408_/B _350_/B 0.13fF
C7754 _501_/a_481_47# _531_/C 0.14fF
C7755 _544_/A _570_/A 0.05fF
C7756 _353_/X _455_/X 0.53fF
C7757 B[1] _417_/A 0.23fF
C7758 VPWR _593_/A 4.79fF
C7759 _586_/a_76_199# _590_/A 0.09fF
C7760 _455_/a_79_199# _542_/D 0.15fF
C7761 _375_/a_222_93# _376_/X 0.00fF
C7762 _445_/A _445_/a_68_297# 0.35fF
C7763 VPWR _542_/A 8.43fF
C7764 _448_/B _324_/a_381_47# 0.02fF
C7765 _544_/A _542_/C 0.27fF
C7766 _480_/Y _486_/X 0.13fF
C7767 _329_/a_226_297# _417_/A 0.02fF
C7768 _538_/A _410_/C 0.04fF
C7769 _573_/Y _593_/Y 0.33fF
C7770 VPWR input4/a_27_47# 0.56fF
C7771 _613_/a_539_297# VPWR 0.02fF
C7772 _411_/B VPWR 0.51fF
C7773 _385_/a_381_47# _393_/A 0.12fF
C7774 _562_/a_493_297# _627_/B 0.08fF
C7775 input12/a_558_47# _442_/D 0.11fF
C7776 input3/a_558_47# VPWR 0.25fF
C7777 _605_/a_80_21# _556_/A 0.10fF
C7778 _497_/A _427_/A 0.00fF
C7779 _528_/a_299_297# _531_/B 0.03fF
C7780 _551_/a_489_413# VPWR 0.39fF
C7781 _633_/Y _585_/B 0.03fF
C7782 _625_/Y _613_/a_227_47# 0.04fF
C7783 _448_/B _378_/A 0.34fF
C7784 _469_/A _469_/X 0.14fF
C7785 _579_/a_145_75# _579_/X 0.02fF
C7786 _436_/A _349_/a_78_199# 0.25fF
C7787 _613_/X _621_/a_78_199# 0.43fF
C7788 _506_/A _442_/A 0.01fF
C7789 _410_/B _455_/X 0.25fF
C7790 _455_/X _456_/a_226_47# 0.52fF
C7791 _381_/C _485_/a_109_47# 0.04fF
C7792 _546_/X _574_/a_299_297# 0.13fF
C7793 _318_/a_197_47# _410_/C 0.03fF
C7794 _516_/A _486_/X 0.60fF
C7795 _519_/X _561_/A 0.15fF
C7796 _539_/A _486_/X 1.67fF
C7797 _367_/a_27_297# _366_/a_76_199# 0.01fF
C7798 _502_/a_493_297# VPWR 0.05fF
C7799 _536_/Y _537_/a_77_199# 0.27fF
C7800 _410_/B _509_/A 0.12fF
C7801 _375_/X _350_/B 0.03fF
C7802 _563_/a_205_297# _542_/D 0.01fF
C7803 _542_/C _391_/B 0.04fF
C7804 _566_/Y _570_/A 0.05fF
C7805 _516_/A _386_/a_558_47# 0.07fF
C7806 A[6] _547_/a_222_93# 0.09fF
C7807 _427_/Y _426_/B 0.31fF
C7808 _512_/a_292_297# VPWR 0.01fF
C7809 _516_/A _513_/A 0.51fF
C7810 _463_/a_489_413# _496_/a_78_199# 0.01fF
C7811 _562_/a_78_199# _627_/C 0.45fF
C7812 _417_/A _383_/X 0.03fF
C7813 _387_/a_215_47# _313_/A 0.22fF
C7814 _569_/A _613_/X 0.05fF
C7815 _576_/a_226_47# _574_/X 0.31fF
C7816 _576_/a_489_413# _575_/X 0.23fF
C7817 _386_/X _518_/a_346_47# 0.02fF
C7818 _396_/X _423_/X 0.10fF
C7819 _458_/X _458_/a_215_47# 0.01fF
C7820 _544_/A _419_/X 0.13fF
C7821 VPWR _366_/a_226_47# 0.08fF
C7822 _545_/a_109_297# _545_/Y 0.02fF
C7823 _353_/X _452_/A 0.09fF
C7824 _544_/A _413_/X 0.06fF
C7825 _611_/X output24/a_27_47# 0.01fF
C7826 B[0] _541_/a_215_47# 0.11fF
C7827 _407_/a_27_47# _406_/B 0.15fF
C7828 _455_/X _376_/X 0.26fF
C7829 _437_/a_79_199# _437_/a_222_93# 0.51fF
C7830 _491_/a_489_413# _489_/X 0.07fF
C7831 _513_/A _478_/a_303_47# 0.03fF
C7832 _520_/X _522_/a_226_297# 0.03fF
C7833 _516_/A _454_/X 0.12fF
C7834 _583_/X M[0] 0.05fF
C7835 _454_/X _539_/A 0.03fF
C7836 _543_/B _588_/A 0.24fF
C7837 _386_/A _479_/a_68_297# 0.02fF
C7838 _566_/A _543_/B 0.17fF
C7839 _631_/B _367_/a_27_297# 0.13fF
C7840 _567_/B _567_/Y 0.50fF
C7841 _570_/B _627_/A 0.26fF
C7842 _613_/X _627_/D 0.80fF
C7843 _567_/B B[0] 0.05fF
C7844 A[6] _518_/X 0.22fF
C7845 _404_/a_664_47# VPWR 0.49fF
C7846 _497_/B VPWR 1.33fF
C7847 _419_/X _391_/B 0.03fF
C7848 _474_/Y _438_/X 0.00fF
C7849 _483_/a_346_47# _410_/C 0.08fF
C7850 _404_/a_558_47# _544_/a_841_47# 0.01fF
C7851 input8/a_27_47# _376_/X 0.01fF
C7852 _375_/X _384_/a_556_47# 0.02fF
C7853 _569_/Y _571_/a_93_21# 0.18fF
C7854 _432_/X _428_/X 0.24fF
C7855 _596_/a_226_47# _601_/A 0.00fF
C7856 _566_/A _565_/a_209_297# 0.04fF
C7857 _627_/X _628_/Y 0.17fF
C7858 A[7] _542_/D 0.06fF
C7859 _563_/a_277_297# _627_/C 0.01fF
C7860 _469_/A _546_/X 0.03fF
C7861 _607_/a_215_47# _618_/A 0.12fF
C7862 _627_/D _609_/a_80_21# 0.24fF
C7863 B[2] input3/a_62_47# 0.01fF
C7864 _626_/Y _548_/X 0.06fF
C7865 _520_/X _483_/X 1.32fF
C7866 _429_/a_76_199# _363_/B 0.17fF
C7867 _381_/C _453_/a_346_47# 0.06fF
C7868 _633_/Y _572_/B 1.04fF
C7869 _417_/a_27_47# _447_/B 0.10fF
C7870 _584_/A _475_/A 0.16fF
C7871 _527_/B _557_/Y 0.01fF
C7872 _595_/a_77_199# _595_/X 0.22fF
C7873 _318_/a_27_47# _318_/a_109_47# 0.03fF
C7874 _327_/a_215_47# _481_/A 0.10fF
C7875 _623_/X _623_/a_76_199# 0.28fF
C7876 _328_/B _336_/a_78_199# 0.00fF
C7877 _530_/a_76_199# VPWR 0.58fF
C7878 VPWR _337_/X 0.96fF
C7879 _376_/X _452_/A 0.69fF
C7880 _567_/B _492_/X 0.24fF
C7881 _500_/a_215_47# _465_/X 0.12fF
C7882 _469_/a_558_47# _469_/a_841_47# 0.07fF
C7883 M[4] _629_/B 0.03fF
C7884 _497_/B _496_/a_215_47# 0.01fF
C7885 _563_/A _381_/B 0.39fF
C7886 _459_/a_76_199# _459_/a_226_47# 0.49fF
C7887 _533_/X _633_/Y 0.03fF
C7888 _611_/a_27_297# _588_/A 0.07fF
C7889 _479_/A _486_/X 0.20fF
C7890 _527_/B _467_/Y 0.38fF
C7891 M[2] _329_/a_76_199# 0.10fF
C7892 _630_/X VPWR 1.38fF
C7893 _340_/A _486_/X 0.56fF
C7894 _587_/A _472_/B 0.78fF
C7895 _456_/a_76_199# _490_/a_78_199# 0.01fF
C7896 _468_/X _436_/X 0.39fF
C7897 _543_/Y _585_/B 0.28fF
C7898 _554_/X _605_/a_80_21# 0.00fF
C7899 _523_/a_226_47# VPWR 0.06fF
C7900 _391_/A _350_/C 0.22fF
C7901 _603_/a_109_297# VPWR 0.01fF
C7902 _513_/A _340_/A 0.07fF
C7903 _542_/a_27_47# _514_/B 0.00fF
C7904 _627_/A _381_/B 0.79fF
C7905 _519_/X VPWR 1.28fF
C7906 _587_/A _436_/a_68_297# 0.30fF
C7907 _488_/a_489_413# VPWR 0.39fF
C7908 _330_/A _406_/A 0.02fF
C7909 _586_/a_76_199# _503_/A 0.22fF
C7910 _360_/X _519_/A 0.03fF
C7911 B[1] _631_/B 0.53fF
C7912 _520_/X A[6] 0.17fF
C7913 _562_/a_493_297# VPWR 0.01fF
C7914 _363_/A _344_/a_78_199# 0.21fF
C7915 _488_/a_226_47# _469_/A 0.07fF
C7916 _525_/a_226_47# _525_/X 0.05fF
C7917 _525_/a_76_199# _524_/X 0.26fF
C7918 _608_/a_215_47# _627_/D 0.07fF
C7919 _352_/a_79_199# _352_/a_448_47# 0.13fF
C7920 _381_/a_27_47# _442_/A 0.22fF
C7921 _390_/B _410_/C 0.54fF
C7922 _476_/a_250_297# _633_/Y 0.21fF
C7923 _351_/X B[5] 0.29fF
C7924 input6/a_27_47# _361_/a_489_413# 0.02fF
C7925 _382_/B _359_/A 0.08fF
C7926 _444_/A _542_/C 0.63fF
C7927 _352_/X _363_/A 0.03fF
C7928 _598_/a_68_297# _597_/a_215_47# 0.01fF
C7929 _536_/Y VPWR 0.51fF
C7930 _386_/a_841_47# _515_/Y 0.04fF
C7931 _423_/a_78_199# _396_/a_93_21# 0.01fF
C7932 _388_/a_27_47# _442_/B 0.54fF
C7933 _542_/B _388_/a_27_47# 0.24fF
C7934 _481_/A _322_/a_27_47# 0.43fF
C7935 _340_/A _454_/X 1.81fF
C7936 _513_/A _566_/A 1.38fF
C7937 _416_/a_78_199# _452_/A 0.50fF
C7938 _586_/a_218_47# _588_/A 0.02fF
C7939 _386_/A _475_/A 0.42fF
C7940 _455_/a_448_47# VPWR 0.03fF
C7941 _581_/B output17/a_27_47# 0.01fF
C7942 _613_/a_77_199# _613_/a_539_297# 0.06fF
C7943 _615_/a_78_199# _616_/B 0.21fF
C7944 _420_/a_222_93# VPWR 0.14fF
C7945 input3/a_62_47# input3/a_381_47# 0.08fF
C7946 _487_/a_292_297# _449_/A 0.01fF
C7947 _432_/a_68_297# _430_/X 0.00fF
C7948 _386_/a_62_47# _386_/A 0.54fF
C7949 _469_/a_381_47# _586_/S 0.04fF
C7950 VPWR _363_/B 2.41fF
C7951 _555_/a_215_297# _554_/B 0.25fF
C7952 _452_/A M[9] 0.07fF
C7953 _551_/a_76_199# _551_/a_226_47# 0.49fF
C7954 _378_/a_558_47# _378_/a_841_47# 0.07fF
C7955 _607_/X _620_/X 0.03fF
C7956 _417_/D _403_/a_27_47# 0.09fF
C7957 _521_/X _488_/X 0.01fF
C7958 _451_/A _340_/A 0.52fF
C7959 _383_/X _631_/B 0.13fF
C7960 _457_/a_489_413# _456_/X 0.16fF
C7961 VPWR _548_/a_226_47# 0.07fF
C7962 _558_/a_77_199# _558_/a_323_297# 0.05fF
C7963 _379_/a_215_47# _542_/D 0.08fF
C7964 _478_/a_27_47# _478_/A 0.44fF
C7965 _483_/a_250_297# _483_/X 0.03fF
C7966 _627_/C _633_/Y 0.03fF
C7967 _445_/X _390_/B 1.03fF
C7968 _626_/Y _523_/X 0.69fF
C7969 _322_/A A[6] 0.06fF
C7970 _349_/a_215_47# VPWR 0.08fF
C7971 _510_/A _503_/A 0.49fF
C7972 _487_/a_215_47# _542_/A 0.02fF
C7973 _538_/Y _559_/X 0.37fF
C7974 _511_/X _522_/a_226_47# 0.09fF
C7975 _522_/X _522_/a_76_199# 0.44fF
C7976 _584_/A _390_/B 0.03fF
C7977 _563_/A _542_/A 0.10fF
C7978 _328_/X _352_/X 0.00fF
C7979 _533_/X _510_/a_68_297# 0.01fF
C7980 _502_/a_78_199# _502_/a_292_297# 0.03fF
C7981 B[7] _598_/A 1.07fF
C7982 _580_/B _579_/a_59_75# 0.37fF
C7983 _500_/a_78_199# _466_/X 0.25fF
C7984 _543_/A _572_/A 0.57fF
C7985 _583_/X _580_/A 0.79fF
C7986 _408_/B _387_/a_215_47# 0.02fF
C7987 _627_/A _542_/A 0.08fF
C7988 _469_/a_664_47# _610_/A 0.10fF
C7989 _411_/B _470_/a_80_21# 0.05fF
C7990 _587_/A _594_/X 0.01fF
C7991 _503_/A _485_/D 0.12fF
C7992 _574_/X _485_/D 0.87fF
C7993 _483_/a_93_21# _483_/a_346_47# 0.05fF
C7994 A[3] _442_/A 1.52fF
C7995 _611_/a_109_297# _633_/Y 0.03fF
C7996 _613_/a_227_47# _586_/S 0.13fF
C7997 VPWR _340_/a_27_47# 0.54fF
C7998 _487_/X _519_/C 0.42fF
C7999 _633_/Y _472_/a_109_297# 0.02fF
C8000 _375_/X _329_/a_226_47# 0.03fF
C8001 _352_/X _374_/X 0.40fF
C8002 _386_/X _475_/A 0.03fF
C8003 _454_/a_76_199# _447_/X 0.44fF
C8004 A[6] _483_/a_250_297# 0.01fF
C8005 input5/a_664_47# _390_/B 0.12fF
C8006 _579_/X _581_/a_27_93# 0.27fF
C8007 M[8] _427_/Y 0.01fF
C8008 _379_/a_493_297# _448_/B 0.02fF
C8009 input6/a_27_47# _361_/a_76_199# 0.00fF
C8010 _485_/D _606_/A 0.15fF
C8011 _632_/a_78_199# _367_/C 0.35fF
C8012 _360_/a_226_47# _360_/a_489_413# 0.02fF
C8013 _360_/a_76_199# _360_/a_226_297# 0.01fF
C8014 _386_/a_62_47# _386_/X 0.41fF
C8015 _344_/a_78_199# _329_/X 0.01fF
C8016 _458_/a_493_297# VPWR 0.01fF
C8017 _410_/B _510_/X 0.56fF
C8018 _410_/B _511_/a_93_21# 0.18fF
C8019 _544_/A _568_/a_227_47# 0.02fF
C8020 _503_/A _483_/X 0.03fF
C8021 _547_/X _469_/X 0.12fF
C8022 _543_/A _542_/D 0.03fF
C8023 _573_/Y _595_/X 0.30fF
C8024 _452_/X _453_/a_250_297# 0.36fF
C8025 _544_/A _382_/A 0.01fF
C8026 _448_/B _519_/A 0.39fF
C8027 _530_/a_226_47# _529_/a_27_47# 0.02fF
C8028 _542_/C _482_/X 0.03fF
C8029 _487_/X _539_/X 0.40fF
C8030 _436_/A _363_/A 0.10fF
C8031 _590_/B _591_/A 0.31fF
C8032 _442_/D _622_/C 0.02fF
C8033 _436_/A _420_/X 0.03fF
C8034 _359_/B _447_/B 0.02fF
C8035 _381_/C _519_/C 1.37fF
C8036 _563_/B _454_/a_76_199# 0.31fF
C8037 _491_/X _525_/a_76_199# 0.01fF
C8038 _476_/X _525_/a_226_47# 0.01fF
C8039 _580_/A _580_/a_68_297# 0.30fF
C8040 _386_/A _390_/B 0.29fF
C8041 _410_/B _443_/a_68_297# 0.07fF
C8042 _386_/X _483_/a_346_47# 0.02fF
C8043 _511_/X _521_/X 0.33fF
C8044 _575_/a_78_199# _540_/X 0.30fF
C8045 _610_/A A[3] 0.03fF
C8046 _597_/a_292_297# _576_/X 0.01fF
C8047 _597_/a_78_199# _575_/X 0.13fF
C8048 _510_/A _471_/Y 1.17fF
C8049 _527_/B _504_/X 0.29fF
C8050 _480_/Y VPWR 1.28fF
C8051 _470_/a_80_21# _470_/a_303_47# 0.04fF
C8052 _415_/a_27_47# _448_/A 0.47fF
C8053 _378_/A _378_/a_62_47# 0.79fF
C8054 _567_/B _456_/X 0.53fF
C8055 _626_/Y _600_/a_27_297# 0.02fF
C8056 VPWR _328_/a_68_297# 0.30fF
C8057 _430_/a_68_297# _430_/X 0.27fF
C8058 VPWR _462_/a_226_47# 0.16fF
C8059 _585_/B _572_/B 0.16fF
C8060 _519_/X _484_/a_292_297# 0.08fF
C8061 _342_/a_68_297# _351_/A 0.00fF
C8062 _417_/D _486_/A 0.21fF
C8063 _583_/X B[0] 0.03fF
C8064 _465_/a_109_297# _427_/Y 0.05fF
C8065 _568_/a_227_47# _566_/Y 0.07fF
C8066 A[6] _503_/A 0.05fF
C8067 _561_/A _340_/A 0.93fF
C8068 _435_/a_27_47# VPWR 0.53fF
C8069 _607_/X VPWR 1.50fF
C8070 _567_/B _478_/A 0.03fF
C8071 _516_/A VPWR 5.48fF
C8072 _390_/D _417_/D 0.74fF
C8073 _360_/X _454_/X 0.02fF
C8074 _544_/A _485_/D 0.44fF
C8075 _442_/B _350_/C 1.61fF
C8076 _328_/B _352_/a_79_199# 0.00fF
C8077 _330_/A _380_/A 3.05fF
C8078 VPWR _539_/A 7.52fF
C8079 _569_/A _571_/a_250_297# 0.03fF
C8080 _363_/A _350_/X 0.62fF
C8081 _360_/a_226_297# _353_/X 0.02fF
C8082 _420_/X _350_/X 0.03fF
C8083 _493_/a_78_199# _460_/a_226_47# 0.00fF
C8084 _510_/A _391_/B 0.03fF
C8085 _347_/A _390_/D 0.03fF
C8086 _404_/a_381_47# _404_/a_558_47# 0.32fF
C8087 VPWR _598_/A 1.23fF
C8088 _510_/A _504_/X 0.40fF
C8089 _539_/X _570_/A 0.03fF
C8090 _587_/A _446_/X 0.18fF
C8091 _626_/a_109_47# _620_/X 0.20fF
C8092 _611_/a_27_297# _592_/a_113_297# 0.02fF
C8093 _382_/X _383_/a_489_413# 0.16fF
C8094 _529_/Y _529_/a_27_47# 0.37fF
C8095 VPWR _489_/X 2.17fF
C8096 _607_/X _606_/Y 0.01fF
C8097 _398_/X B[5] 0.04fF
C8098 B[7] _588_/A 0.84fF
C8099 _314_/X _328_/a_68_297# 0.21fF
C8100 _366_/a_226_47# _368_/A 0.05fF
C8101 _534_/a_303_47# _485_/D 0.03fF
C8102 _386_/A _471_/A 0.02fF
C8103 _616_/Y _625_/a_27_297# 0.02fF
C8104 _563_/B _447_/X 0.44fF
C8105 _383_/a_226_297# _452_/A 0.02fF
C8106 _492_/a_226_47# _524_/X 0.01fF
C8107 _442_/B _367_/C 0.09fF
C8108 _424_/X _422_/X 0.08fF
C8109 _330_/A _384_/a_226_47# 0.02fF
C8110 _542_/B _442_/A 0.03fF
C8111 _470_/a_209_297# _411_/X 0.02fF
C8112 _332_/a_68_297# _332_/X 0.27fF
C8113 _547_/X _546_/X 3.80fF
C8114 _550_/a_215_47# _511_/X 0.03fF
C8115 _442_/B _442_/A 0.63fF
C8116 _386_/X _390_/B 0.07fF
C8117 _574_/X _598_/B 0.12fF
C8118 _563_/D _406_/A 0.13fF
C8119 _437_/a_79_199# _437_/X 0.29fF
C8120 _519_/X _563_/A 0.00fF
C8121 _566_/Y _485_/D 0.17fF
C8122 _572_/a_68_297# VPWR 0.41fF
C8123 _532_/a_76_199# VPWR 0.57fF
C8124 _368_/B _337_/A 0.03fF
C8125 _487_/X _381_/C 0.48fF
C8126 _509_/Y _511_/a_584_47# 0.01fF
C8127 M[12] input12/a_558_47# 0.07fF
C8128 _578_/a_78_199# _578_/a_292_297# 0.03fF
C8129 _588_/A _574_/a_81_21# 0.12fF
C8130 _417_/D _324_/a_62_47# 0.23fF
C8131 _328_/A _332_/X 0.03fF
C8132 _519_/A _314_/a_68_297# 0.33fF
C8133 _554_/A _555_/a_298_297# 0.11fF
C8134 _503_/A _609_/a_209_47# 0.01fF
C8135 _534_/a_80_21# _386_/a_558_47# 0.00fF
C8136 _368_/a_68_297# _368_/a_150_297# 0.02fF
C8137 _554_/X _556_/A 0.29fF
C8138 _433_/Y _472_/B 1.77fF
C8139 _488_/a_489_413# _627_/A 0.09fF
C8140 _568_/a_77_199# VPWR 0.89fF
C8141 _570_/a_68_297# _570_/a_150_297# 0.02fF
C8142 _360_/X _337_/A 0.03fF
C8143 _590_/A _590_/B 2.90fF
C8144 _427_/Y _428_/X 0.02fF
C8145 _544_/A A[6] 0.03fF
C8146 _561_/A _454_/a_489_413# 0.00fF
C8147 _540_/a_250_297# _535_/Y 0.00fF
C8148 _432_/a_68_297# _430_/a_68_297# 0.02fF
C8149 _490_/X _446_/X 0.17fF
C8150 _533_/a_77_199# _533_/a_539_297# 0.06fF
C8151 _455_/X _382_/B 0.27fF
C8152 _487_/X _570_/A 0.41fF
C8153 _412_/X _458_/a_78_199# 0.35fF
C8154 _426_/B _427_/A 0.07fF
C8155 _449_/A _628_/Y 0.01fF
C8156 _390_/D _445_/a_150_297# 0.01fF
C8157 _629_/A VPWR 1.79fF
C8158 _443_/A _390_/a_27_47# 0.00fF
C8159 _567_/B _493_/a_78_199# 0.18fF
C8160 _609_/a_80_21# _609_/a_303_47# 0.04fF
C8161 _410_/B _511_/X 0.01fF
C8162 _627_/C _585_/B 0.32fF
C8163 _542_/C _487_/X 0.03fF
C8164 _368_/A _337_/X 0.28fF
C8165 _350_/X _374_/X 0.16fF
C8166 _618_/A _624_/X 0.01fF
C8167 _421_/a_76_199# _421_/a_489_413# 0.12fF
C8168 _611_/X _622_/C 0.10fF
C8169 _563_/D _350_/C 0.40fF
C8170 _386_/X _471_/A 0.39fF
C8171 _623_/X _584_/A 0.27fF
C8172 _530_/X _486_/X 0.08fF
C8173 _410_/B _390_/B 1.35fF
C8174 B[3] VPWR 0.45fF
C8175 _397_/X _399_/a_78_199# 0.34fF
C8176 _594_/a_27_297# _593_/A 0.20fF
C8177 _479_/A VPWR 0.36fF
C8178 _324_/a_664_47# _324_/a_841_47# 0.29fF
C8179 _340_/A VPWR 3.86fF
C8180 _417_/A _633_/Y 0.03fF
C8181 _583_/X _625_/a_27_47# 0.08fF
C8182 _612_/A _588_/Y 2.01fF
C8183 _513_/A _530_/X 0.09fF
C8184 _625_/Y _442_/D 0.03fF
C8185 _474_/Y _510_/A 0.31fF
C8186 _380_/A _442_/B 0.03fF
C8187 _611_/a_27_297# _611_/a_373_47# 0.08fF
C8188 _499_/a_81_21# _497_/A 0.17fF
C8189 _353_/a_68_297# _445_/A 0.33fF
C8190 _472_/Y _503_/A 0.09fF
C8191 _628_/a_28_47# _572_/A 0.01fF
C8192 _578_/a_215_47# _549_/X 0.14fF
C8193 _452_/X _449_/A 1.83fF
C8194 _487_/X _535_/A 0.02fF
C8195 _563_/A _349_/a_215_47# 0.11fF
C8196 input5/a_381_47# VPWR 0.30fF
C8197 _365_/a_81_21# _630_/a_76_199# 0.00fF
C8198 _583_/X _616_/A 0.27fF
C8199 _444_/Y _445_/X 0.02fF
C8200 _588_/A VPWR 4.77fF
C8201 _530_/X _486_/a_150_297# 0.02fF
C8202 M[5] _397_/X 0.04fF
C8203 _502_/a_215_47# _494_/X 0.05fF
C8204 _563_/D _442_/A 0.03fF
C8205 _600_/a_27_297# _593_/A 0.13fF
C8206 _386_/X _446_/a_256_47# 0.03fF
C8207 _452_/A _378_/a_558_47# 0.17fF
C8208 _599_/A _598_/a_68_297# 0.27fF
C8209 _544_/a_664_47# _588_/A 0.05fF
C8210 _549_/a_76_199# _549_/a_226_47# 0.49fF
C8211 _362_/a_226_47# _363_/B 0.05fF
C8212 _390_/a_27_47# _390_/a_109_47# 0.03fF
C8213 _566_/A VPWR 3.77fF
C8214 _625_/Y _588_/Y 1.94fF
C8215 _424_/X _478_/A 0.06fF
C8216 _599_/A _599_/Y 0.35fF
C8217 _557_/A _602_/Y 0.26fF
C8218 _454_/X _530_/X 0.21fF
C8219 _567_/Y _469_/A 0.03fF
C8220 _627_/C _447_/X 0.01fF
C8221 _567_/B _570_/B 0.08fF
C8222 B[7] _559_/X 0.03fF
C8223 _626_/a_109_47# VPWR 0.23fF
C8224 _488_/a_76_199# _488_/a_226_47# 0.49fF
C8225 _424_/a_226_47# _424_/a_489_413# 0.02fF
C8226 _424_/a_76_199# _424_/a_226_297# 0.01fF
C8227 _567_/B _626_/Y 0.03fF
C8228 _542_/C _570_/A 0.10fF
C8229 _403_/a_27_47# _410_/C 0.10fF
C8230 _382_/B _452_/A 0.88fF
C8231 _602_/A _581_/B 0.06fF
C8232 _548_/a_226_47# _548_/X 0.05fF
C8233 _548_/a_76_199# _547_/X 0.49fF
C8234 _391_/B _391_/a_68_297# 0.30fF
C8235 B[0] _469_/A 0.60fF
C8236 _443_/A _391_/B 0.01fF
C8237 _562_/a_78_199# _562_/a_292_297# 0.03fF
C8238 _620_/X _616_/B 0.23fF
C8239 _347_/A _563_/a_27_297# 0.01fF
C8240 VPWR _521_/a_493_297# 0.01fF
C8241 _618_/Y _618_/A 0.59fF
C8242 _626_/a_397_297# _623_/X 0.22fF
C8243 _543_/B _514_/B 0.64fF
C8244 _330_/A B[4] 0.24fF
C8245 _476_/X _492_/a_489_413# 0.16fF
C8246 _491_/X _492_/a_226_47# 0.54fF
C8247 _426_/A _350_/X 0.19fF
C8248 _622_/a_29_53# _622_/X 0.20fF
C8249 _622_/a_111_297# _627_/B 0.02fF
C8250 _544_/A _418_/B 0.50fF
C8251 _533_/a_539_297# _469_/X 0.08fF
C8252 _410_/B _471_/A 0.05fF
C8253 _570_/X _503_/A 0.36fF
C8254 _536_/Y _537_/a_227_47# 0.15fF
C8255 _569_/A A[3] 1.00fF
C8256 _627_/C _563_/B 1.57fF
C8257 VPWR _398_/a_76_199# 0.43fF
C8258 _608_/a_292_297# _627_/B 0.01fF
C8259 _396_/a_250_297# _631_/B 0.12fF
C8260 _426_/A _478_/A 0.03fF
C8261 B[7] _616_/B 0.92fF
C8262 _565_/a_80_21# _514_/A 0.01fF
C8263 _567_/B _406_/Y 0.18fF
C8264 _476_/a_93_21# _476_/a_256_47# 0.03fF
C8265 _570_/A _535_/A 0.39fF
C8266 M[6] output29/a_27_47# 0.46fF
C8267 _419_/X _421_/a_226_47# 0.31fF
C8268 _630_/a_489_413# _629_/a_68_297# 0.02fF
C8269 _539_/a_68_297# A[3] 0.24fF
C8270 _605_/a_209_297# _557_/Y 0.02fF
C8271 _338_/a_79_199# _366_/a_489_413# 0.03fF
C8272 _338_/a_222_93# _366_/a_226_47# 0.00fF
C8273 _552_/a_76_199# _552_/a_489_413# 0.12fF
C8274 _633_/Y _469_/X 0.10fF
C8275 _458_/X _436_/X 0.79fF
C8276 _540_/a_93_21# _539_/X 0.19fF
C8277 input16/a_27_47# _549_/a_76_199# 0.02fF
C8278 _452_/A _632_/a_78_199# 0.01fF
C8279 _510_/a_68_297# _533_/a_77_199# 0.01fF
C8280 _454_/a_489_413# VPWR 0.17fF
C8281 _523_/a_226_47# _523_/X 0.05fF
C8282 _471_/Y _472_/Y 0.79fF
C8283 _444_/Y _386_/A 0.20fF
C8284 VPWR _344_/a_292_297# 0.02fF
C8285 _603_/a_109_297# _603_/Y 0.02fF
C8286 _437_/X _503_/A 0.24fF
C8287 _443_/A _441_/a_78_199# 0.21fF
C8288 output30/a_27_47# VPWR 0.68fF
C8289 _620_/a_226_297# _618_/Y 0.01fF
C8290 _417_/D _628_/Y 0.08fF
C8291 _455_/a_79_199# _455_/a_448_47# 0.13fF
C8292 _485_/A _334_/a_303_47# 0.09fF
C8293 VPWR _558_/a_539_297# 0.02fF
C8294 VPWR _554_/a_68_297# 0.33fF
C8295 _627_/D A[3] 0.03fF
C8296 _594_/X _540_/X 0.01fF
C8297 _567_/B _381_/B 0.40fF
C8298 _487_/X _477_/a_493_297# 0.02fF
C8299 _510_/A _387_/a_78_199# 0.18fF
C8300 _375_/a_448_47# _375_/X 0.01fF
C8301 _455_/X _442_/B 1.01fF
C8302 _542_/B _455_/X 0.03fF
C8303 _583_/X M[11] 0.25fF
C8304 _370_/A _337_/X 0.01fF
C8305 _416_/a_78_199# _418_/A 0.31fF
C8306 _538_/A _535_/Y 0.37fF
C8307 _336_/a_78_199# _328_/A 0.17fF
C8308 _581_/B _606_/A 0.07fF
C8309 _510_/A _385_/a_841_47# 0.05fF
C8310 _516_/A _563_/A 0.12fF
C8311 _611_/X _612_/A 0.19fF
C8312 _623_/a_76_199# _628_/Y 0.05fF
C8313 _567_/B _527_/A 0.88fF
C8314 M[8] _467_/Y 0.38fF
C8315 _503_/A _439_/a_76_199# 0.03fF
C8316 _572_/A _574_/a_299_297# 0.12fF
C8317 _418_/A M[9] 0.25fF
C8318 _417_/D _452_/X 0.03fF
C8319 _612_/Y _624_/a_76_199# 0.05fF
C8320 _435_/a_27_47# _627_/A 0.07fF
C8321 _368_/B VPWR 1.56fF
C8322 _583_/X _619_/Y 0.19fF
C8323 _448_/A _453_/a_256_47# 0.03fF
C8324 _577_/a_226_47# _390_/D 0.07fF
C8325 _627_/A _539_/A 0.51fF
C8326 _559_/X VPWR 2.52fF
C8327 VPWR _550_/a_292_297# 0.01fF
C8328 _493_/a_493_297# _458_/X 0.08fF
C8329 _338_/a_222_93# _337_/X 0.13fF
C8330 _611_/X _625_/Y 0.72fF
C8331 _613_/X _623_/X 1.12fF
C8332 _417_/D _481_/a_27_47# 0.09fF
C8333 _446_/a_93_21# _446_/a_250_297# 0.50fF
C8334 _615_/a_292_297# _593_/A 0.02fF
C8335 _513_/A _514_/B 0.14fF
C8336 _351_/A _408_/B 0.38fF
C8337 _369_/a_76_199# _369_/a_489_413# 0.12fF
C8338 _360_/X VPWR 4.88fF
C8339 _612_/A _618_/A 0.20fF
C8340 VPWR _625_/a_277_47# 0.04fF
C8341 _605_/a_209_297# _606_/A 0.04fF
C8342 _610_/A _591_/A 0.95fF
C8343 _506_/Y _503_/A 0.20fF
C8344 _448_/B _561_/A 0.82fF
C8345 _413_/X _419_/X 0.19fF
C8346 _557_/A _558_/X 1.26fF
C8347 _608_/X _627_/C 0.10fF
C8348 _421_/a_76_199# _421_/X 0.22fF
C8349 _446_/X _433_/Y 0.03fF
C8350 _469_/a_558_47# _545_/Y 0.08fF
C8351 _523_/a_226_297# _631_/Y 0.01fF
C8352 B[4] _442_/B 0.13fF
C8353 _390_/D _410_/C 2.02fF
C8354 _444_/Y _386_/X 1.60fF
C8355 _633_/Y _546_/X 0.12fF
C8356 _385_/a_664_47# _475_/A 0.12fF
C8357 VPWR _465_/X 2.10fF
C8358 _485_/A _542_/D 0.19fF
C8359 _504_/X _525_/X 1.38fF
C8360 _633_/Y _631_/B 0.03fF
C8361 VPWR _409_/a_215_47# 0.05fF
C8362 _475_/X _478_/A 0.08fF
C8363 VPWR _616_/B 2.92fF
C8364 _342_/X _344_/a_292_297# 0.01fF
C8365 _349_/a_78_199# _349_/a_215_47# 0.26fF
C8366 _493_/a_215_47# _493_/X 0.01fF
C8367 _586_/S _564_/a_219_297# 0.19fF
C8368 _444_/A _443_/A 0.24fF
C8369 _610_/A _624_/a_206_369# 0.04fF
C8370 VPWR _571_/a_93_21# 0.37fF
C8371 _625_/Y _618_/A 0.01fF
C8372 _566_/Y _570_/X 0.85fF
C8373 _503_/A _559_/a_77_199# 0.43fF
C8374 _429_/a_226_47# _350_/X 0.31fF
C8375 B[7] _530_/X 0.03fF
C8376 _396_/a_93_21# _396_/a_346_47# 0.05fF
C8377 _567_/B _542_/A 0.03fF
C8378 M[8] _427_/A 0.15fF
C8379 _601_/Y _618_/A 0.34fF
C8380 _599_/A _616_/A 0.15fF
C8381 _613_/a_77_199# _588_/A 0.30fF
C8382 _568_/a_227_297# _433_/Y 0.04fF
C8383 _347_/A _355_/A 0.19fF
C8384 _633_/Y _411_/X 0.12fF
C8385 _455_/X _563_/D 0.03fF
C8386 _469_/A _572_/A 0.26fF
C8387 _527_/B _556_/A 0.13fF
C8388 _451_/A _514_/B 0.03fF
C8389 _375_/X _351_/A 0.18fF
C8390 _352_/X _383_/X 0.08fF
C8391 _424_/X _406_/Y 0.06fF
C8392 _416_/a_78_199# _416_/a_215_47# 0.26fF
C8393 _328_/A _410_/C 0.02fF
C8394 _611_/a_109_297# _627_/C 0.02fF
C8395 _587_/A _592_/a_199_47# 0.02fF
C8396 _608_/a_292_297# VPWR 0.01fF
C8397 _550_/X VPWR 1.73fF
C8398 _584_/A _486_/A 0.21fF
C8399 _480_/Y _505_/a_209_297# 0.09fF
C8400 _519_/C _485_/D 0.03fF
C8401 _449_/A _447_/B 0.16fF
C8402 _520_/X _442_/A 0.18fF
C8403 _620_/a_489_413# VPWR 0.39fF
C8404 _391_/A _475_/A 0.00fF
C8405 _390_/D _445_/X 1.01fF
C8406 _465_/X _501_/Y 0.97fF
C8407 _380_/A _518_/X 0.03fF
C8408 _474_/Y _472_/Y 0.10fF
C8409 _416_/a_215_47# M[9] 0.12fF
C8410 _390_/D _584_/A 0.03fF
C8411 _563_/A _340_/A 0.04fF
C8412 _442_/D _433_/Y 0.05fF
C8413 _482_/a_68_297# _481_/A 0.08fF
C8414 _544_/A _544_/a_62_47# 0.52fF
C8415 VPWR _592_/a_113_297# 0.59fF
C8416 _444_/Y _410_/B 0.85fF
C8417 VPWR M[10] 0.92fF
C8418 _538_/A A[3] 0.22fF
C8419 _388_/a_27_47# _390_/a_27_47# 0.01fF
C8420 _586_/S _442_/D 0.03fF
C8421 _448_/a_68_297# _453_/a_250_297# 0.03fF
C8422 _634_/Y _369_/a_489_413# 0.00fF
C8423 _627_/X _625_/Y 0.25fF
C8424 _505_/a_303_47# _481_/A 0.03fF
C8425 _360_/X _342_/X 0.16fF
C8426 _534_/a_80_21# VPWR 0.32fF
C8427 A[6] _482_/X 0.11fF
C8428 _565_/a_80_21# _512_/a_215_47# 0.00fF
C8429 _417_/D _479_/a_150_297# 0.02fF
C8430 _465_/a_109_297# _427_/A 0.04fF
C8431 _504_/a_227_47# _468_/a_215_47# 0.07fF
C8432 _331_/a_27_47# _384_/a_226_47# 0.02fF
C8433 _539_/A _508_/a_227_47# 0.02fF
C8434 _411_/B _411_/A 0.50fF
C8435 _417_/A _447_/X 0.18fF
C8436 _389_/a_27_47# _410_/C 0.00fF
C8437 _425_/a_489_413# _478_/A 0.09fF
C8438 _623_/a_76_199# _623_/a_226_297# 0.01fF
C8439 _432_/A _371_/a_68_297# 0.33fF
C8440 VPWR _553_/a_215_47# 0.07fF
C8441 _627_/A _588_/A 0.94fF
C8442 _441_/a_78_199# _441_/a_292_297# 0.03fF
C8443 _563_/D _477_/a_215_47# 0.13fF
C8444 A[5] _398_/X 0.05fF
C8445 _436_/A B[1] 1.75fF
C8446 _338_/X _419_/X 0.26fF
C8447 _466_/a_78_199# _466_/X 0.21fF
C8448 _583_/X _626_/Y 0.02fF
C8449 B[2] _616_/Y 0.12fF
C8450 _566_/A _627_/A 0.27fF
C8451 B[0] M[6] 0.03fF
C8452 _404_/a_62_47# _588_/A 0.02fF
C8453 _539_/X _483_/X 0.52fF
C8454 _594_/a_27_297# _594_/a_373_47# 0.08fF
C8455 _585_/B _469_/X 0.48fF
C8456 _502_/a_78_199# _492_/X 0.01fF
C8457 _587_/A _436_/X 0.34fF
C8458 _458_/a_78_199# _458_/a_292_297# 0.03fF
C8459 _431_/a_76_199# VPWR 0.49fF
C8460 _410_/C _316_/a_558_47# 0.24fF
C8461 _448_/B VPWR 5.23fF
C8462 _610_/A _590_/A 1.59fF
C8463 _404_/a_664_47# _543_/A 0.07fF
C8464 _408_/B _519_/A 1.09fF
C8465 _497_/B _567_/B 0.12fF
C8466 _588_/A _548_/X 0.01fF
C8467 _347_/A _313_/a_27_47# 0.02fF
C8468 _500_/a_78_199# _498_/A 0.03fF
C8469 _322_/A _442_/A 0.34fF
C8470 _442_/D _442_/a_27_47# 0.28fF
C8471 _523_/X _489_/X 0.02fF
C8472 A[6] _519_/C 0.12fF
C8473 _406_/A _503_/A 0.27fF
C8474 _386_/A _390_/D 0.03fF
C8475 _543_/Y _546_/X 0.22fF
C8476 _444_/A _446_/a_250_297# 0.21fF
C8477 _567_/Y _547_/X 0.48fF
C8478 VPWR _530_/X 10.63fF
C8479 _343_/a_226_47# _343_/X 0.21fF
C8480 _565_/a_80_21# _417_/D 0.11fF
C8481 _591_/Y _590_/B 0.05fF
C8482 _380_/A _520_/X 0.03fF
C8483 _476_/X _504_/X 0.37fF
C8484 B[0] _547_/X 0.03fF
C8485 _533_/X _533_/a_77_199# 0.22fF
C8486 _347_/A _565_/a_80_21# 0.12fF
C8487 _433_/a_109_297# VPWR 0.01fF
C8488 _422_/a_226_47# _421_/X 0.55fF
C8489 _599_/A _619_/Y 0.22fF
C8490 _487_/X _485_/D 0.42fF
C8491 _567_/Y _570_/a_68_297# 0.08fF
C8492 _510_/A _438_/X 0.66fF
C8493 _373_/a_113_297# _373_/Y 0.42fF
C8494 _614_/a_226_47# _612_/Y 0.07fF
C8495 _440_/X _458_/X 2.32fF
C8496 _576_/a_76_199# _576_/a_489_413# 0.12fF
C8497 _422_/X _407_/Y 0.03fF
C8498 B[2] _620_/a_76_199# 0.11fF
C8499 A[6] _539_/X 0.08fF
C8500 _350_/a_27_297# _442_/B 0.05fF
C8501 _429_/a_76_199# input14/a_27_47# 0.01fF
C8502 _632_/a_78_199# _475_/A 0.38fF
C8503 _432_/A _432_/X 0.03fF
C8504 _436_/A _383_/X 0.74fF
C8505 B[1] _350_/X 0.94fF
C8506 _390_/B _432_/X 0.03fF
C8507 _439_/X _503_/A 0.02fF
C8508 _328_/A _352_/a_79_199# 0.29fF
C8509 _392_/A _350_/B 0.05fF
C8510 _562_/a_215_47# _564_/A 0.01fF
C8511 _373_/a_113_297# VPWR 0.55fF
C8512 _621_/a_78_199# _591_/A 0.25fF
C8513 _375_/X _519_/A 2.24fF
C8514 _531_/A _558_/X 0.03fF
C8515 _474_/A _587_/A 0.34fF
C8516 _519_/a_29_53# _447_/B 0.01fF
C8517 _376_/X _356_/a_78_199# 0.03fF
C8518 _383_/X _542_/D 0.39fF
C8519 _633_/a_74_47# _632_/a_78_199# 0.00fF
C8520 _573_/A _590_/B 0.01fF
C8521 _381_/C _485_/D 0.15fF
C8522 _417_/D _447_/B 0.04fF
C8523 _318_/a_27_47# _380_/A 0.02fF
C8524 _424_/a_226_47# _406_/A 0.01fF
C8525 _424_/a_76_199# _406_/B 0.01fF
C8526 _487_/X _483_/X 0.32fF
C8527 _465_/X _531_/C 0.01fF
C8528 _380_/A _384_/a_489_413# 0.09fF
C8529 _563_/B _484_/a_215_47# 0.10fF
C8530 _605_/a_80_21# _605_/a_209_297# 0.16fF
C8531 _397_/a_76_199# _397_/X 0.24fF
C8532 _507_/Y _472_/B 0.03fF
C8533 _499_/a_299_297# _467_/Y 0.18fF
C8534 _363_/A _630_/X 0.13fF
C8535 _513_/a_27_47# _542_/a_27_47# 0.05fF
C8536 _442_/D _316_/a_664_47# 0.29fF
C8537 _358_/a_197_47# _442_/A 0.12fF
C8538 _442_/D _443_/B 0.16fF
C8539 B[0] _488_/a_76_199# 0.09fF
C8540 _423_/a_292_297# VPWR 0.01fF
C8541 _585_/B _546_/X 0.09fF
C8542 _493_/a_292_297# VPWR 0.01fF
C8543 _322_/A _380_/A 0.29fF
C8544 _614_/a_76_199# _610_/Y 0.10fF
C8545 _627_/D _586_/a_505_21# 0.01fF
C8546 _367_/a_27_297# _367_/a_205_297# 0.01fF
C8547 _604_/X _604_/a_209_297# 0.11fF
C8548 _423_/a_215_47# _384_/X 0.03fF
C8549 _485_/D _570_/A 1.91fF
C8550 _567_/B _536_/Y 0.00fF
C8551 _386_/X _390_/D 0.75fF
C8552 VPWR _557_/B 2.02fF
C8553 _383_/X _350_/X 0.03fF
C8554 _384_/a_489_413# _384_/a_226_47# 0.02fF
C8555 _600_/a_27_297# _598_/A 0.21fF
C8556 _342_/X _369_/a_226_297# 0.01fF
C8557 _572_/B _469_/X 0.03fF
C8558 output21/a_27_47# _583_/X 0.19fF
C8559 _362_/a_489_413# _352_/X 0.02fF
C8560 VPWR _453_/a_93_21# 0.39fF
C8561 _527_/B _497_/A 0.08fF
C8562 _542_/C _485_/D 0.03fF
C8563 _382_/A _419_/X 0.07fF
C8564 _503_/A _442_/A 0.03fF
C8565 _487_/X A[6] 0.13fF
C8566 _631_/Y _410_/C 1.68fF
C8567 _613_/X _612_/Y 0.44fF
C8568 _509_/Y _533_/a_77_199# 0.17fF
C8569 _469_/a_558_47# _622_/C 0.09fF
C8570 output20/a_27_47# _607_/X 0.63fF
C8571 _390_/D _575_/X 0.04fF
C8572 _524_/a_493_297# VPWR 0.01fF
C8573 _314_/a_68_297# VPWR 0.25fF
C8574 _538_/Y _472_/B 0.56fF
C8575 M[2] _343_/X 0.23fF
C8576 _547_/a_222_93# _547_/a_448_47# 0.03fF
C8577 _516_/a_27_47# _516_/A 0.32fF
C8578 _627_/D _591_/A 1.60fF
C8579 _418_/X _378_/a_381_47# 0.17fF
C8580 _533_/X _551_/a_226_47# 0.06fF
C8581 VPWR input14/a_27_47# 0.52fF
C8582 _551_/X _551_/a_76_199# 0.37fF
C8583 _474_/Y _476_/X 0.11fF
C8584 _563_/A _409_/a_215_47# 0.16fF
C8585 A[2] _606_/A 0.08fF
C8586 M[10] _531_/C 0.00fF
C8587 _406_/A _391_/B 0.13fF
C8588 _420_/a_222_93# _420_/X 0.05fF
C8589 _475_/A _442_/B 0.07fF
C8590 _559_/X _548_/X 1.21fF
C8591 _631_/A _384_/a_76_199# 0.04fF
C8592 _363_/A _363_/B 1.00fF
C8593 _510_/A _419_/X 0.02fF
C8594 _381_/C A[6] 1.51fF
C8595 _485_/D _535_/A 1.06fF
C8596 _448_/a_68_297# _449_/A 0.27fF
C8597 _440_/a_226_297# _436_/X 0.01fF
C8598 _556_/Y VPWR 1.43fF
C8599 _488_/a_226_47# _585_/B 0.01fF
C8600 _513_/a_303_47# _542_/C 0.06fF
C8601 _481_/a_27_47# _410_/C 0.07fF
C8602 _503_/a_558_47# _446_/X 0.08fF
C8603 _361_/a_226_47# _361_/X 0.13fF
C8604 _476_/a_250_297# _469_/X 0.03fF
C8605 _615_/a_78_199# _594_/X 0.34fF
C8606 _368_/B _368_/A 2.51fF
C8607 _407_/Y _478_/A 0.18fF
C8608 _583_/X _542_/A 0.22fF
C8609 _627_/A _571_/a_93_21# 0.11fF
C8610 _360_/X _362_/a_226_47# 0.02fF
C8611 _524_/a_215_47# _490_/X 0.10fF
C8612 _314_/a_68_297# _314_/X 0.27fF
C8613 _485_/A _381_/B 0.94fF
C8614 _584_/A _628_/Y 0.17fF
C8615 _469_/A _570_/B 0.34fF
C8616 _381_/C _358_/a_303_47# 0.03fF
C8617 _626_/Y _469_/A 0.03fF
C8618 _611_/X _610_/Y 0.06fF
C8619 _315_/a_161_47# _563_/B 0.33fF
C8620 _630_/X _374_/X 0.88fF
C8621 _410_/B _390_/D 1.97fF
C8622 _371_/a_68_297# _371_/A 0.33fF
C8623 _445_/X _631_/Y 0.03fF
C8624 _610_/A _503_/A 0.10fF
C8625 _518_/X _547_/a_448_47# 0.22fF
C8626 _488_/a_226_297# _486_/X 0.01fF
C8627 _342_/a_68_297# VPWR 0.33fF
C8628 _583_/X input3/a_558_47# 0.10fF
C8629 VPWR _514_/B 1.21fF
C8630 A[6] _570_/A 0.09fF
C8631 _520_/a_226_47# _547_/a_79_199# 0.00fF
C8632 _486_/X _472_/B 0.50fF
C8633 _360_/a_489_413# _375_/a_79_199# 0.01fF
C8634 _431_/a_556_47# _430_/X 0.02fF
C8635 _431_/a_226_297# _428_/X 0.02fF
C8636 VPWR _467_/a_109_297# 0.01fF
C8637 _624_/a_76_199# _624_/a_489_47# 0.14fF
C8638 _623_/a_226_47# _621_/X 0.31fF
C8639 _404_/a_381_47# _572_/A 0.14fF
C8640 _595_/a_227_47# _469_/X 0.01fF
C8641 _542_/C A[6] 0.05fF
C8642 _383_/a_226_47# VPWR 0.10fF
C8643 output19/a_27_47# M[15] 0.28fF
C8644 M[11] output23/a_27_47# 0.02fF
C8645 _544_/A _367_/C 0.05fF
C8646 M[8] _465_/a_27_297# 0.20fF
C8647 _608_/a_493_297# _586_/S 0.02fF
C8648 _610_/A _609_/a_209_297# 0.04fF
C8649 _462_/X VPWR 1.79fF
C8650 _572_/B _546_/X 0.33fF
C8651 _546_/a_76_199# _544_/a_381_47# 0.01fF
C8652 _382_/X _420_/a_544_297# 0.04fF
C8653 _608_/X _469_/X 0.06fF
C8654 _516_/A _379_/a_215_47# 0.10fF
C8655 _514_/a_68_297# _514_/A 0.32fF
C8656 _355_/A _410_/C 0.03fF
C8657 _457_/a_226_47# _446_/X 0.25fF
C8658 _423_/a_78_199# _383_/X 0.13fF
C8659 _382_/X _420_/a_79_199# 0.18fF
C8660 _627_/X _433_/Y 0.05fF
C8661 _420_/a_448_47# _452_/A 0.09fF
C8662 _385_/a_381_47# VPWR 0.31fF
C8663 _480_/A _479_/B 0.02fF
C8664 _509_/Y _469_/X 0.97fF
C8665 _419_/X _631_/A 1.53fF
C8666 _610_/Y _618_/A 0.12fF
C8667 _523_/X _554_/a_68_297# 0.20fF
C8668 _627_/X _586_/S 0.07fF
C8669 _569_/A _590_/A 0.07fF
C8670 _454_/X _472_/B 0.03fF
C8671 _337_/B _519_/A 0.58fF
C8672 _549_/X _540_/X 0.03fF
C8673 _412_/a_76_199# VPWR 0.50fF
C8674 _520_/a_76_199# _518_/X 0.39fF
C8675 _467_/a_109_297# _501_/Y 0.02fF
C8676 _371_/A _432_/X 0.11fF
C8677 _570_/X _539_/X 0.00fF
C8678 _629_/B _430_/X 0.38fF
C8679 _420_/X _458_/a_493_297# 0.08fF
C8680 _510_/A _336_/a_493_297# 0.09fF
C8681 _469_/A _381_/B 0.08fF
C8682 _394_/a_558_47# _394_/a_664_47# 0.60fF
C8683 _394_/a_381_47# _394_/a_841_47# 0.03fF
C8684 _407_/a_109_297# VPWR 0.01fF
C8685 _417_/D _418_/X 0.33fF
C8686 _479_/B _481_/A 0.18fF
C8687 _464_/Y _466_/X 0.17fF
C8688 _496_/a_493_297# _461_/X 0.08fF
C8689 _496_/a_215_47# _462_/X 0.05fF
C8690 _563_/D _475_/A 0.03fF
C8691 B[0] _480_/A 0.46fF
C8692 _386_/A _631_/Y 0.03fF
C8693 _562_/a_215_47# _451_/A 0.01fF
C8694 _630_/X _426_/A 1.31fF
C8695 _465_/a_27_297# _465_/a_109_297# 0.45fF
C8696 _628_/a_382_297# _623_/a_76_199# 0.05fF
C8697 _347_/A _445_/A 0.26fF
C8698 _445_/A _332_/X 0.01fF
C8699 _590_/A _627_/D 0.95fF
C8700 _569_/Y _588_/Y 0.16fF
C8701 _576_/a_226_47# _485_/D 0.07fF
C8702 _390_/B _442_/B 0.29fF
C8703 _485_/a_27_47# _486_/A 0.10fF
C8704 _542_/B _390_/B 0.47fF
C8705 _610_/A _590_/a_150_297# 0.02fF
C8706 _313_/A VPWR 1.58fF
C8707 _563_/A _530_/X 0.05fF
C8708 _410_/B _389_/a_27_47# 0.12fF
C8709 _410_/a_109_47# VPWR 0.01fF
C8710 _411_/a_68_297# _386_/X 0.14fF
C8711 _342_/a_68_297# _342_/X 0.27fF
C8712 _485_/A _542_/A 0.19fF
C8713 _408_/B _337_/A 0.06fF
C8714 _420_/X _328_/a_68_297# 0.07fF
C8715 _469_/a_381_47# VPWR 0.35fF
C8716 _567_/Y _633_/Y 0.07fF
C8717 B[0] _481_/A 0.66fF
C8718 _335_/a_62_47# _510_/A 0.47fF
C8719 _627_/A _530_/X 0.03fF
C8720 _439_/X _474_/Y 0.02fF
C8721 _564_/a_219_297# _564_/A 0.22fF
C8722 _469_/a_62_47# _469_/A 0.44fF
C8723 B[0] _633_/Y 0.05fF
C8724 _473_/a_323_297# _472_/B 0.11fF
C8725 _385_/a_664_47# _394_/a_841_47# 0.02fF
C8726 _393_/A _394_/a_62_47# 0.00fF
C8727 _544_/A _380_/A 0.34fF
C8728 _390_/a_197_47# _442_/B 0.03fF
C8729 _315_/a_161_47# _627_/C 0.03fF
C8730 _542_/C _390_/a_109_47# 0.02fF
C8731 _343_/a_76_199# VPWR 0.57fF
C8732 _633_/Y _521_/a_292_297# 0.08fF
C8733 _368_/B _370_/A 0.03fF
C8734 _546_/a_76_199# _546_/a_226_297# 0.01fF
C8735 _546_/a_226_47# _546_/a_489_413# 0.02fF
C8736 _455_/X _503_/A 0.12fF
C8737 _520_/a_76_199# _520_/X 0.22fF
C8738 _387_/a_78_199# _387_/a_292_297# 0.03fF
C8739 _530_/X _548_/X 0.12fF
C8740 _383_/a_76_199# _383_/X 0.22fF
C8741 _489_/a_226_47# _488_/X 0.50fF
C8742 _489_/a_489_413# _483_/X 0.25fF
C8743 _426_/A _363_/B 0.01fF
C8744 _501_/a_397_297# _531_/A 0.12fF
C8745 _378_/a_62_47# VPWR 0.53fF
C8746 _527_/B _532_/a_489_47# 0.02fF
C8747 _328_/B _442_/B 0.06fF
C8748 _503_/A _509_/A 0.12fF
C8749 _567_/B _532_/a_76_199# 0.05fF
C8750 _614_/a_226_47# output24/a_27_47# 0.01fF
C8751 _375_/X _337_/A 0.03fF
C8752 _483_/a_93_21# _481_/a_27_47# 0.00fF
C8753 _440_/a_76_199# _440_/a_226_47# 0.49fF
C8754 _455_/a_222_93# _542_/D 0.02fF
C8755 _328_/X _328_/a_68_297# 0.28fF
C8756 _557_/A _531_/A 0.78fF
C8757 _386_/X _631_/Y 0.07fF
C8758 _567_/B _460_/a_556_47# 0.02fF
C8759 _386_/A _355_/A 0.03fF
C8760 _629_/B _432_/a_68_297# 0.05fF
C8761 _517_/a_68_297# VPWR 0.31fF
C8762 _417_/a_27_47# _519_/A 0.26fF
C8763 _613_/a_227_47# VPWR 0.09fF
C8764 _419_/X _418_/B 0.00fF
C8765 _383_/X _381_/B 0.48fF
C8766 _385_/a_558_47# _393_/A 0.24fF
C8767 _562_/a_215_47# _627_/B 0.10fF
C8768 input12/a_664_47# _442_/D 0.05fF
C8769 input3/a_664_47# VPWR 0.37fF
C8770 _510_/a_68_297# _510_/a_150_297# 0.02fF
C8771 _568_/a_77_199# _567_/B 0.50fF
C8772 _413_/X _418_/B 0.02fF
C8773 _413_/a_68_297# _413_/a_150_297# 0.02fF
C8774 _623_/X A[3] 0.05fF
C8775 _563_/B _452_/a_68_297# 0.34fF
C8776 _311_/a_27_47# _447_/B 0.40fF
C8777 _537_/a_77_199# _472_/B 0.35fF
C8778 _614_/a_556_47# _591_/A 0.02fF
C8779 _533_/X M[0] 0.10fF
C8780 _436_/A _349_/a_292_297# 0.02fF
C8781 _407_/Y _406_/Y 0.79fF
C8782 output26/a_27_47# B[5] 0.11fF
C8783 _541_/a_215_47# _340_/A 0.19fF
C8784 _455_/X _456_/a_489_413# 0.14fF
C8785 _390_/D _506_/A 0.48fF
C8786 _563_/D _390_/B 0.09fF
C8787 _542_/C _446_/a_250_297# 0.00fF
C8788 _584_/A _313_/a_27_47# 0.10fF
C8789 _591_/Y _610_/A 0.19fF
C8790 _466_/a_78_199# _431_/X 0.42fF
C8791 VPWR _575_/a_78_199# 0.62fF
C8792 _437_/X _438_/X 1.17fF
C8793 _367_/a_27_297# _366_/a_226_47# 0.03fF
C8794 _502_/a_215_47# VPWR 0.13fF
C8795 _563_/a_277_297# _542_/D 0.01fF
C8796 _570_/X _570_/A 0.25fF
C8797 _512_/a_493_297# VPWR 0.01fF
C8798 _516_/A _386_/a_664_47# 0.12fF
C8799 _386_/X _481_/a_27_47# 0.22fF
C8800 _329_/a_76_199# _343_/a_489_413# 0.02fF
C8801 _559_/a_77_199# _539_/X 0.38fF
C8802 _516_/A _355_/a_161_47# 0.60fF
C8803 _543_/B _442_/D 0.03fF
C8804 _517_/X _486_/X 0.09fF
C8805 _355_/A _483_/a_93_21# 0.01fF
C8806 _629_/A _363_/A 0.14fF
C8807 _448_/B _419_/a_489_413# 0.01fF
C8808 _427_/Y _390_/B 0.61fF
C8809 input1/a_27_47# A[0] 0.32fF
C8810 M[2] _371_/B 0.24fF
C8811 _444_/A _442_/A 0.41fF
C8812 _630_/a_226_47# _371_/A 0.00fF
C8813 _630_/a_489_413# _629_/B 0.00fF
C8814 _503_/a_62_47# _503_/A 0.51fF
C8815 _543_/A _340_/A 0.03fF
C8816 _569_/A _503_/A 0.31fF
C8817 _455_/X _471_/Y 0.09fF
C8818 _347_/A _441_/a_215_47# 0.12fF
C8819 _576_/a_489_413# _574_/X 0.07fF
C8820 _523_/X _553_/a_215_47# 0.11fF
C8821 _600_/a_27_297# _616_/B 0.02fF
C8822 _542_/A _489_/a_76_199# 0.02fF
C8823 _603_/Y _553_/a_215_47# 0.02fF
C8824 VPWR _366_/a_489_413# 0.39fF
C8825 _545_/Y _584_/A 1.12fF
C8826 _544_/A _455_/X 0.75fF
C8827 _613_/X output24/a_27_47# 0.09fF
C8828 _491_/a_226_297# _489_/X 0.05fF
C8829 _417_/D _587_/A 0.05fF
C8830 _538_/A _520_/X 0.57fF
C8831 _439_/a_76_199# _438_/X 0.30fF
C8832 _350_/X _432_/B 0.03fF
C8833 _440_/a_76_199# _439_/X 0.21fF
C8834 _597_/a_215_47# _598_/A 0.01fF
C8835 _410_/B _631_/Y 0.64fF
C8836 _567_/B _588_/A 0.53fF
C8837 _387_/a_78_199# _350_/C 0.36fF
C8838 _529_/a_27_47# _531_/B 0.01fF
C8839 _567_/B _566_/A 0.49fF
C8840 _584_/A _326_/A 0.03fF
C8841 _386_/X _355_/A 0.40fF
C8842 _543_/Y B[0] 0.03fF
C8843 B[0] _515_/Y 0.10fF
C8844 _627_/D _503_/A 0.09fF
C8845 _519_/X _485_/A 0.65fF
C8846 _603_/Y _530_/X 0.03fF
C8847 _607_/a_493_297# _606_/A 0.04fF
C8848 _607_/a_78_199# _601_/A 0.40fF
C8849 _430_/X _428_/X 2.24fF
C8850 _567_/Y _521_/a_78_199# 0.01fF
C8851 _382_/B _356_/a_78_199# 0.18fF
C8852 _367_/a_27_297# _337_/X 0.01fF
C8853 B[0] _521_/a_78_199# 0.04fF
C8854 _487_/X _559_/a_77_199# 0.12fF
C8855 _533_/a_77_199# _469_/X 0.18fF
C8856 _446_/X _454_/X 0.03fF
C8857 _570_/B _547_/X 0.17fF
C8858 _627_/D _609_/a_209_297# 0.14fF
C8859 _615_/a_215_47# _585_/B 0.30fF
C8860 _554_/X _581_/B 0.03fF
C8861 _547_/a_79_199# _486_/B 0.27fF
C8862 _591_/A _601_/A 0.04fF
C8863 _565_/a_80_21# _386_/A 0.14fF
C8864 _533_/X _533_/a_227_47# 0.04fF
C8865 _520_/X _488_/X 0.13fF
C8866 _429_/a_226_47# _363_/B 0.06fF
C8867 _521_/a_78_199# _521_/a_292_297# 0.03fF
C8868 _633_/Y _572_/A 0.90fF
C8869 _625_/Y _623_/a_76_199# 0.01fF
C8870 _536_/a_109_297# _587_/A 0.02fF
C8871 _376_/X _382_/X 2.82fF
C8872 _386_/a_62_47# _520_/X 0.10fF
C8873 _502_/a_78_199# _527_/A 0.21fF
C8874 _544_/A _477_/a_215_47# 0.33fF
C8875 _570_/B _570_/a_68_297# 0.30fF
C8876 _390_/D _535_/Y 0.56fF
C8877 _503_/a_62_47# _471_/Y 0.16fF
C8878 _500_/a_215_47# _466_/X 0.18fF
C8879 _544_/A _452_/A 0.24fF
C8880 _530_/a_226_47# VPWR 0.14fF
C8881 _457_/X _460_/X 0.07fF
C8882 _469_/a_664_47# _469_/a_841_47# 0.29fF
C8883 _442_/D _486_/X 0.03fF
C8884 _380_/A B[5] 0.04fF
C8885 _459_/a_76_199# _459_/a_489_413# 0.12fF
C8886 _624_/a_76_199# _624_/X 0.23fF
C8887 _408_/B VPWR 4.17fF
C8888 _544_/A _569_/A 0.44fF
C8889 _548_/a_489_413# _574_/a_81_21# 0.02fF
C8890 _456_/a_226_47# _490_/a_78_199# 0.01fF
C8891 _506_/Y _508_/a_77_199# 0.17fF
C8892 _337_/B _337_/A 0.33fF
C8893 _510_/A _631_/A 0.66fF
C8894 _386_/a_664_47# _479_/A 0.00fF
C8895 _523_/a_489_413# VPWR 0.39fF
C8896 _567_/Y _585_/B 0.15fF
C8897 _584_/A _486_/a_68_297# 0.02fF
C8898 _355_/a_161_47# _340_/A 0.15fF
C8899 _330_/A A[0] 0.02fF
C8900 B[0] _585_/B 0.62fF
C8901 _513_/A _417_/a_27_47# 0.29fF
C8902 _562_/a_215_47# VPWR 0.05fF
C8903 VPWR _472_/B 4.20fF
C8904 _352_/a_222_93# _352_/a_448_47# 0.03fF
C8905 _488_/a_489_413# _469_/A 0.02fF
C8906 _525_/a_226_47# _524_/X 0.55fF
C8907 input6/a_27_47# VPWR 0.54fF
C8908 _559_/a_77_199# _570_/A 0.22fF
C8909 _563_/A _313_/A 0.03fF
C8910 _480_/A _478_/A 0.00fF
C8911 _433_/Y _431_/X 0.21fF
C8912 _603_/Y _557_/B 0.04fF
C8913 VPWR _445_/a_68_297# 0.28fF
C8914 _454_/X _442_/D 0.48fF
C8915 _607_/X _583_/X 0.27fF
C8916 _381_/B _547_/X 0.10fF
C8917 _544_/A _547_/a_448_47# 0.16fF
C8918 VPWR _436_/a_68_297# 0.27fF
C8919 _459_/X _460_/X 0.11fF
C8920 _408_/B _314_/X 0.35fF
C8921 _560_/a_27_47# _381_/C 0.01fF
C8922 _569_/A _566_/Y 0.93fF
C8923 _359_/B _519_/A 0.03fF
C8924 _456_/X _633_/Y 0.72fF
C8925 _579_/a_59_75# _606_/A 0.30fF
C8926 _353_/a_68_297# _519_/A 0.43fF
C8927 _596_/a_76_199# B[7] 0.01fF
C8928 _521_/a_215_47# _486_/X 0.11fF
C8929 _400_/a_80_21# _392_/Y 0.23fF
C8930 _611_/a_27_297# _614_/a_76_199# 0.00fF
C8931 _469_/a_558_47# _433_/Y 0.15fF
C8932 _554_/X _476_/X 0.00fF
C8933 _402_/a_27_47# _438_/X 0.00fF
C8934 _613_/a_77_199# _613_/a_227_47# 0.24fF
C8935 _583_/a_76_199# _582_/Y 0.25fF
C8936 VPWR output22/a_27_47# 0.64fF
C8937 _375_/X VPWR 4.68fF
C8938 _445_/A _410_/C 0.33fF
C8939 _487_/a_78_199# _519_/C 0.12fF
C8940 _487_/a_493_297# _449_/A 0.01fF
C8941 _381_/B _570_/a_68_297# 0.08fF
C8942 _509_/Y _533_/a_227_47# 0.05fF
C8943 input3/a_62_47# input3/a_558_47# 0.03fF
C8944 _567_/B _559_/X 0.58fF
C8945 _454_/a_76_199# _454_/a_226_47# 0.49fF
C8946 _386_/a_381_47# _386_/A 0.15fF
C8947 _629_/B _629_/a_68_297# 0.35fF
C8948 _469_/a_558_47# _586_/S 0.02fF
C8949 _329_/a_76_199# _442_/B 0.02fF
C8950 _555_/a_298_297# _554_/B 0.24fF
C8951 _529_/Y VPWR 0.76fF
C8952 _580_/A _533_/X 0.42fF
C8953 _378_/a_664_47# _378_/a_841_47# 0.29fF
C8954 _629_/A _426_/A 0.05fF
C8955 A[6] _485_/D 1.22fF
C8956 _551_/a_76_199# _551_/a_489_413# 0.12fF
C8957 _633_/Y _478_/A 0.03fF
C8958 _347_/A _387_/a_215_47# 0.11fF
C8959 _417_/A _631_/B 0.31fF
C8960 _456_/X _490_/a_215_47# 0.07fF
C8961 VPWR _554_/A 1.37fF
C8962 _616_/Y _599_/Y 0.58fF
C8963 _520_/X _511_/X 0.15fF
C8964 _513_/a_27_47# _513_/A 0.65fF
C8965 _516_/A output32/a_27_47# 0.01fF
C8966 output30/a_27_47# _558_/a_77_199# 0.03fF
C8967 _544_/A _379_/a_78_199# 0.32fF
C8968 _448_/a_68_297# _311_/a_27_47# 0.00fF
C8969 VPWR _548_/a_489_413# 0.39fF
C8970 _558_/a_77_199# _558_/a_539_297# 0.06fF
C8971 _603_/Y _556_/Y 0.17fF
C8972 _398_/a_76_199# _374_/X 0.45fF
C8973 _564_/a_219_297# _627_/B 0.09fF
C8974 _360_/X _363_/A 0.03fF
C8975 _538_/A _503_/A 0.32fF
C8976 _488_/a_76_199# _381_/B 0.10fF
C8977 A[6] _483_/X 0.11fF
C8978 _444_/A _455_/X 0.80fF
C8979 _375_/X _314_/X 1.07fF
C8980 _522_/X _522_/a_226_47# 0.24fF
C8981 _510_/X _503_/A 0.28fF
C8982 _360_/X _420_/X 0.03fF
C8983 _503_/A _511_/a_93_21# 0.01fF
C8984 _529_/a_27_47# _498_/A 0.03fF
C8985 _442_/A _539_/X 0.15fF
C8986 _563_/A _517_/a_68_297# 0.20fF
C8987 _567_/B _571_/a_93_21# 0.03fF
C8988 _412_/X _631_/B 0.45fF
C8989 _635_/a_27_413# B[5] 0.07fF
C8990 _423_/a_78_199# _396_/X 0.39fF
C8991 _543_/Y _572_/A 0.08fF
C8992 _411_/B _470_/a_209_297# 0.06fF
C8993 _519_/a_29_53# _484_/a_78_199# 0.01fF
C8994 _445_/A _445_/X 0.05fF
C8995 _587_/A _595_/X 0.01fF
C8996 B[1] _363_/B 0.07fF
C8997 _417_/D _484_/a_78_199# 0.18fF
C8998 _612_/Y A[3] 0.03fF
C8999 _445_/A _584_/A 0.19fF
C9000 _390_/D A[3] 0.05fF
C9001 _611_/a_27_297# _611_/X 0.34fF
C9002 _613_/a_227_47# _627_/A 0.16fF
C9003 _513_/A _358_/a_27_47# 0.15fF
C9004 input5/a_841_47# _390_/B 0.07fF
C9005 _454_/a_76_199# _453_/X 0.24fF
C9006 _454_/a_226_47# _447_/X 0.25fF
C9007 _584_/A _395_/a_68_297# 0.35fF
C9008 _591_/Y _627_/D 0.60fF
C9009 _318_/a_27_47# _390_/B 0.02fF
C9010 M[7] _557_/Y 0.78fF
C9011 _439_/X _438_/X 0.63fF
C9012 _379_/a_215_47# _448_/B 0.15fF
C9013 _542_/A _547_/X 0.12fF
C9014 _594_/X VPWR 1.90fF
C9015 _344_/a_215_47# _343_/X 0.17fF
C9016 _412_/X _411_/X 0.01fF
C9017 _516_/A _485_/A 0.30fF
C9018 _386_/a_381_47# _386_/X 0.71fF
C9019 _584_/A _622_/C 0.30fF
C9020 _458_/a_215_47# VPWR 0.07fF
C9021 _411_/A _409_/a_215_47# 0.01fF
C9022 _587_/a_27_47# _627_/D 0.22fF
C9023 _375_/X _342_/X 0.03fF
C9024 _410_/B _511_/a_250_297# 0.04fF
C9025 _499_/a_81_21# _499_/a_299_297# 0.21fF
C9026 _543_/Y _542_/D 0.01fF
C9027 _546_/X _469_/X 0.27fF
C9028 _467_/Y M[7] 0.04fF
C9029 _487_/a_78_199# _487_/X 0.21fF
C9030 _442_/D _627_/B 0.92fF
C9031 _590_/B _621_/X 0.02fF
C9032 _378_/a_381_47# _324_/a_381_47# 0.01fF
C9033 A[5] _399_/a_78_199# 0.02fF
C9034 _596_/a_76_199# VPWR 0.51fF
C9035 _563_/B _454_/a_226_47# 0.02fF
C9036 _490_/X _525_/a_76_199# 0.01fF
C9037 _491_/X _525_/a_226_47# 0.01fF
C9038 _443_/a_68_297# _390_/a_27_47# 0.01fF
C9039 _410_/B _443_/a_150_297# 0.01fF
C9040 _585_/B _616_/A 0.01fF
C9041 _510_/a_68_297# _478_/A 0.03fF
C9042 _530_/a_226_47# _531_/C 0.00fF
C9043 _522_/X _521_/X 0.49fF
C9044 _545_/Y _590_/a_68_297# 0.00fF
C9045 _575_/a_78_199# _548_/X 0.42fF
C9046 _510_/X _471_/Y 0.01fF
C9047 _313_/a_27_47# _395_/X 0.00fF
C9048 _510_/A _472_/Y 0.92fF
C9049 _527_/B _525_/X 0.01fF
C9050 _583_/X _588_/A 0.05fF
C9051 _597_/a_493_297# _576_/X 0.01fF
C9052 _597_/a_78_199# _574_/X 0.01fF
C9053 _597_/a_215_47# _559_/X 0.03fF
C9054 _378_/A _378_/a_381_47# 0.02fF
C9055 _442_/D _620_/X 0.05fF
C9056 _632_/a_78_199# _632_/a_215_47# 0.26fF
C9057 _573_/Y _591_/A 0.02fF
C9058 _360_/X _374_/X 1.09fF
C9059 _623_/X _591_/A 0.10fF
C9060 VPWR _462_/a_489_413# 0.42fF
C9061 _585_/B _572_/A 4.08fF
C9062 A[5] M[5] 0.79fF
C9063 _381_/C _367_/C 0.09fF
C9064 _465_/a_109_47# _427_/Y 0.01fF
C9065 _384_/X _397_/X 0.09fF
C9066 _417_/D _433_/Y 0.05fF
C9067 _386_/A _390_/a_303_47# 0.03fF
C9068 B[7] _442_/D 0.03fF
C9069 _513_/A _359_/B 0.21fF
C9070 _406_/A _419_/X 0.09fF
C9071 _447_/X _453_/X 3.21fF
C9072 _554_/X _555_/a_27_413# 0.62fF
C9073 _381_/C _442_/A 1.14fF
C9074 _577_/a_76_199# VPWR 0.51fF
C9075 _328_/B _352_/a_222_93# 0.00fF
C9076 _337_/B VPWR 1.52fF
C9077 _376_/X _447_/B 0.03fF
C9078 _469_/A _539_/A 0.02fF
C9079 _587_/A _410_/C 0.16fF
C9080 _597_/a_215_47# _616_/B 0.27fF
C9081 _625_/a_27_297# _625_/a_27_47# 0.07fF
C9082 _467_/Y _390_/B 0.13fF
C9083 _497_/A _497_/a_68_297# 0.30fF
C9084 _404_/a_381_47# _404_/a_664_47# 0.09fF
C9085 _461_/a_493_297# _390_/B 0.02fF
C9086 VPWR _517_/X 0.75fF
C9087 _567_/B _530_/X 0.09fF
C9088 _626_/a_109_297# _620_/X 0.02fF
C9089 _607_/X _599_/A 0.49fF
C9090 _623_/a_76_199# _433_/Y 0.08fF
C9091 _385_/a_664_47# _631_/Y 0.16fF
C9092 _417_/D _540_/X 0.07fF
C9093 _359_/B _454_/X 0.45fF
C9094 _538_/A _566_/Y 0.01fF
C9095 B[0] _627_/C 0.07fF
C9096 _616_/Y _625_/a_27_47# 0.02fF
C9097 _376_/X _376_/a_68_297# 0.27fF
C9098 _423_/X _422_/X 1.36fF
C9099 _563_/B _453_/X 0.19fF
C9100 _492_/a_489_413# _524_/X 0.01fF
C9101 _443_/a_68_297# _391_/B 0.01fF
C9102 M[5] _629_/a_68_297# 0.08fF
C9103 _599_/A _598_/A 0.03fF
C9104 _378_/A _512_/a_215_47# 0.11fF
C9105 input10/a_27_47# _397_/X 0.01fF
C9106 _529_/Y _531_/C 0.30fF
C9107 _563_/A _408_/B 0.58fF
C9108 _442_/A _508_/a_77_199# 0.08fF
C9109 _456_/a_76_199# _454_/X 0.31fF
C9110 _442_/A _316_/a_62_47# 0.45fF
C9111 _446_/X VPWR 4.49fF
C9112 _503_/A _511_/X 0.05fF
C9113 _542_/C _442_/A 1.77fF
C9114 _550_/a_215_47# _522_/X 0.05fF
C9115 _409_/a_78_199# _409_/a_215_47# 0.26fF
C9116 _390_/D _442_/B 0.03fF
C9117 _564_/a_219_297# VPWR 0.23fF
C9118 _616_/Y _616_/A 0.79fF
C9119 _589_/a_226_47# _588_/Y 0.53fF
C9120 _542_/B _390_/D 0.46fF
C9121 _572_/a_150_297# VPWR 0.00fF
C9122 _437_/a_222_93# _437_/X 0.05fF
C9123 _570_/X _485_/D 0.14fF
C9124 _568_/a_323_297# _587_/A 0.04fF
C9125 _532_/a_206_369# VPWR 0.10fF
C9126 _487_/X _380_/A 2.71fF
C9127 _536_/a_109_297# _433_/Y 0.04fF
C9128 _473_/a_77_199# _503_/A 0.02fF
C9129 _510_/A _437_/X 0.01fF
C9130 M[12] input12/a_664_47# 0.12fF
C9131 _493_/X _459_/X 0.01fF
C9132 _588_/A _574_/a_299_297# 0.18fF
C9133 _562_/a_215_47# _563_/A 0.11fF
C9134 _390_/B _503_/A 0.69fF
C9135 _419_/X _350_/C 0.37fF
C9136 _475_/A _391_/B 0.03fF
C9137 _503_/A _609_/a_303_47# 0.01fF
C9138 _513_/A _534_/a_209_297# 0.01fF
C9139 _633_/Y _385_/a_62_47# 0.10fF
C9140 _442_/B _332_/a_68_297# 0.12fF
C9141 _585_/B _478_/A 0.04fF
C9142 _568_/a_227_297# VPWR 0.01fF
C9143 _587_/A _584_/A 0.06fF
C9144 _631_/B _411_/X 0.60fF
C9145 _584_/A _612_/A 0.02fF
C9146 _519_/a_29_53# _378_/A 0.14fF
C9147 _447_/X _542_/D 0.15fF
C9148 M[9] _447_/B 0.74fF
C9149 _381_/B _481_/A 0.32fF
C9150 _627_/A _472_/B 2.05fF
C9151 _533_/a_77_199# _533_/a_227_47# 0.24fF
C9152 _381_/C _380_/A 1.19fF
C9153 _417_/D _378_/A 1.19fF
C9154 _438_/a_68_297# _472_/B 0.31fF
C9155 _489_/X _489_/a_76_199# 0.22fF
C9156 _606_/A _601_/A 0.45fF
C9157 _419_/X _367_/C 0.05fF
C9158 _572_/B _572_/A 1.24fF
C9159 _328_/A _442_/B 0.54fF
C9160 _390_/B _427_/A 0.17fF
C9161 _519_/X _547_/X 0.00fF
C9162 _347_/A _378_/A 0.14fF
C9163 _567_/B _557_/B 0.08fF
C9164 _545_/a_109_297# VPWR 0.01fF
C9165 _347_/A _346_/a_161_47# 0.68fF
C9166 _353_/a_68_297# _337_/A 0.01fF
C9167 _429_/a_76_199# _398_/a_226_47# 0.01fF
C9168 _429_/a_226_47# _398_/a_76_199# 0.01fF
C9169 _421_/a_226_47# _421_/a_489_413# 0.02fF
C9170 _421_/a_76_199# _421_/a_226_297# 0.01fF
C9171 _353_/X _445_/A 0.02fF
C9172 _613_/X _622_/C 0.32fF
C9173 _399_/a_78_199# _398_/X 0.28fF
C9174 _623_/X _590_/A 0.14fF
C9175 _625_/Y _584_/A 1.31fF
C9176 _595_/a_77_199# _503_/A 0.17fF
C9177 _442_/D VPWR 4.11fF
C9178 _563_/B _542_/D 0.81fF
C9179 _390_/B _390_/a_27_47# 0.56fF
C9180 _594_/a_109_297# _593_/A 0.12fF
C9181 VPWR _522_/a_76_199# 0.45fF
C9182 _579_/X VPWR 1.79fF
C9183 _380_/A _570_/A 0.20fF
C9184 _380_/A _351_/X 0.06fF
C9185 _536_/Y _547_/X 0.10fF
C9186 _380_/A _384_/a_76_199# 0.08fF
C9187 _629_/X _630_/X 0.01fF
C9188 _516_/A _356_/a_215_47# 0.08fF
C9189 _417_/a_27_47# VPWR 0.57fF
C9190 _492_/a_76_199# VPWR 0.52fF
C9191 _498_/Y VPWR 1.90fF
C9192 _628_/a_300_47# _572_/A 0.02fF
C9193 _471_/A _503_/A 0.70fF
C9194 _499_/a_299_297# _497_/A 0.14fF
C9195 _419_/X _632_/a_493_297# 0.04fF
C9196 _578_/a_215_47# _580_/B 0.01fF
C9197 _533_/X _551_/X 2.92fF
C9198 _586_/a_505_21# _469_/a_841_47# 0.01fF
C9199 _609_/a_80_21# _622_/C 0.24fF
C9200 input5/a_558_47# VPWR 0.22fF
C9201 _365_/a_81_21# _630_/a_226_47# 0.02fF
C9202 M[5] _398_/X 0.06fF
C9203 _473_/a_77_199# _471_/Y 0.14fF
C9204 _588_/Y VPWR 3.40fF
C9205 _386_/X _446_/a_346_47# 0.02fF
C9206 _469_/A _588_/A 0.88fF
C9207 _471_/Y _390_/B 0.11fF
C9208 _363_/A input14/a_27_47# 0.14fF
C9209 _620_/a_76_199# _620_/a_226_47# 0.49fF
C9210 _390_/D _563_/D 1.16fF
C9211 _384_/a_76_199# _384_/a_226_47# 0.49fF
C9212 _549_/a_76_199# _549_/a_489_413# 0.12fF
C9213 _382_/B _382_/X 0.28fF
C9214 _611_/X B[7] 0.05fF
C9215 _480_/A _542_/A 0.13fF
C9216 _557_/Y _604_/a_80_21# 0.10fF
C9217 _476_/X _510_/A 0.53fF
C9218 _375_/a_79_199# _375_/a_222_93# 0.51fF
C9219 _566_/A _469_/A 0.03fF
C9220 _628_/Y M[15] 0.04fF
C9221 _626_/a_109_297# VPWR 0.01fF
C9222 _488_/a_76_199# _488_/a_489_413# 0.12fF
C9223 _316_/a_62_47# _316_/a_381_47# 0.08fF
C9224 _548_/a_226_47# _547_/X 0.46fF
C9225 _548_/a_76_199# _546_/X 0.32fF
C9226 _508_/a_77_199# _508_/a_227_297# 0.13fF
C9227 _527_/B _528_/a_81_21# 0.02fF
C9228 _619_/Y _616_/Y 0.14fF
C9229 _543_/B _514_/A 0.34fF
C9230 _620_/X _618_/A 1.48fF
C9231 _543_/A _514_/B 0.10fF
C9232 VPWR _521_/a_215_47# 0.06fF
C9233 _476_/X _492_/a_226_297# 0.01fF
C9234 _491_/X _492_/a_489_413# 0.16fF
C9235 _557_/B _558_/a_77_199# 0.55fF
C9236 _626_/a_397_297# _625_/Y 0.12fF
C9237 _537_/a_227_47# _472_/B 0.11fF
C9238 A[5] _380_/A 0.17fF
C9239 _613_/X _589_/a_76_199# 0.22fF
C9240 _533_/a_227_47# _469_/X 0.03fF
C9241 _533_/X _456_/X 0.03fF
C9242 _544_/A _418_/A 0.11fF
C9243 _444_/A _443_/a_68_297# 0.52fF
C9244 B[2] _580_/A 0.12fF
C9245 _513_/a_27_47# VPWR 0.78fF
C9246 _481_/A _542_/A 0.03fF
C9247 _608_/X _572_/A 0.45fF
C9248 _539_/a_68_297# _539_/X 0.27fF
C9249 VPWR _398_/a_226_47# 0.06fF
C9250 _380_/A _419_/X 0.03fF
C9251 _633_/Y _593_/A 0.09fF
C9252 _506_/Y _483_/X 0.10fF
C9253 _431_/a_76_199# _426_/A 0.07fF
C9254 _390_/B _391_/B 0.02fF
C9255 _455_/X _381_/C 0.03fF
C9256 _608_/a_493_297# _627_/B 0.08fF
C9257 _440_/X _460_/a_76_199# 0.63fF
C9258 _567_/B _462_/X 0.01fF
C9259 _633_/Y _542_/A 0.36fF
C9260 _614_/a_76_199# VPWR 0.46fF
C9261 _476_/a_93_21# _476_/a_346_47# 0.05fF
C9262 _342_/a_68_297# _420_/X 0.07fF
C9263 _627_/B _627_/a_27_297# 0.41fF
C9264 _419_/X _421_/a_489_413# 0.07fF
C9265 _545_/Y _515_/A 0.01fF
C9266 _411_/B _633_/Y 0.13fF
C9267 _533_/X _478_/A 0.03fF
C9268 _590_/a_68_297# _622_/C 0.02fF
C9269 _627_/C _572_/A 1.35fF
C9270 _338_/a_222_93# _366_/a_489_413# 0.01fF
C9271 _540_/a_250_297# _539_/X 0.31fF
C9272 _630_/X _432_/B 0.31fF
C9273 _552_/a_226_47# _552_/a_489_413# 0.02fF
C9274 _552_/a_76_199# _552_/a_226_297# 0.01fF
C9275 _614_/a_226_47# _625_/Y 0.05fF
C9276 _614_/a_489_413# _623_/X 0.06fF
C9277 _612_/Y _586_/a_505_21# 0.00fF
C9278 _608_/a_78_199# _608_/X 0.23fF
C9279 input16/a_27_47# _549_/a_226_47# 0.00fF
C9280 _471_/Y _471_/A 0.57fF
C9281 _545_/Y _546_/a_76_199# 0.28fF
C9282 _627_/X _627_/B 0.14fF
C9283 _349_/a_78_199# _408_/B 0.18fF
C9284 _634_/Y _368_/B 0.13fF
C9285 _430_/a_68_297# _430_/a_150_297# 0.02fF
C9286 VPWR _344_/a_493_297# 0.01fF
C9287 _410_/B _446_/a_346_47# 0.08fF
C9288 input7/a_27_47# VPWR 0.53fF
C9289 _603_/a_27_47# _603_/Y 0.22fF
C9290 _395_/a_68_297# _395_/X 0.27fF
C9291 _455_/a_222_93# _455_/a_448_47# 0.03fF
C9292 _556_/Y _558_/a_77_199# 0.34fF
C9293 VPWR _558_/a_227_47# 0.04fF
C9294 _620_/a_76_199# _619_/Y 0.22fF
C9295 _608_/X _542_/D 0.64fF
C9296 _608_/a_78_199# _627_/C 0.45fF
C9297 _375_/a_79_199# _455_/X 0.17fF
C9298 _335_/a_62_47# _367_/C 0.01fF
C9299 _515_/Y _381_/B 1.43fF
C9300 _461_/a_78_199# VPWR 0.64fF
C9301 _485_/a_27_47# _486_/B 0.19fF
C9302 _553_/a_78_199# _553_/a_215_47# 0.26fF
C9303 _570_/B _585_/B 0.44fF
C9304 _612_/Y _591_/A 0.33fF
C9305 _506_/Y A[6] 0.06fF
C9306 _542_/C _455_/X 0.72fF
C9307 _393_/A _584_/A 0.01fF
C9308 _368_/B _367_/a_27_297# 0.20fF
C9309 _423_/a_78_199# _423_/X 0.21fF
C9310 _627_/C _542_/D 3.28fF
C9311 _416_/a_78_199# _418_/X 0.06fF
C9312 _358_/a_27_47# VPWR 0.79fF
C9313 _508_/a_77_199# _509_/A 0.22fF
C9314 input13/a_27_47# _374_/a_78_199# 0.01fF
C9315 _613_/X _612_/A 0.53fF
C9316 _471_/A _446_/a_93_21# 0.01fF
C9317 _503_/A _439_/a_226_47# 0.08fF
C9318 _595_/a_77_199# _566_/Y 0.28fF
C9319 _572_/A _574_/a_384_47# 0.12fF
C9320 _338_/a_79_199# _332_/X 0.01fF
C9321 _418_/X M[9] 0.05fF
C9322 _627_/X B[7] 0.06fF
C9323 _612_/Y _624_/a_206_369# 0.05fF
C9324 _563_/A _517_/X 0.53fF
C9325 input15/a_75_212# VPWR 0.56fF
C9326 _432_/B _363_/B 0.28fF
C9327 _518_/X _486_/A 0.08fF
C9328 _587_/a_27_47# _601_/A 0.03fF
C9329 _611_/X VPWR 2.19fF
C9330 VPWR _550_/a_493_297# 0.01fF
C9331 _576_/X VPWR 1.07fF
C9332 _493_/a_215_47# _458_/X 0.10fF
C9333 _386_/a_381_47# _515_/A 0.16fF
C9334 _428_/a_81_21# _427_/Y 0.51fF
C9335 _542_/B _631_/Y 1.53fF
C9336 _442_/B _631_/Y 0.48fF
C9337 _613_/X _625_/Y 0.60fF
C9338 _544_/a_381_47# _503_/A 0.00fF
C9339 _513_/A _514_/A 0.01fF
C9340 _375_/X _396_/a_93_21# 0.01fF
C9341 _573_/Y _574_/X 0.16fF
C9342 _446_/a_93_21# _446_/a_256_47# 0.03fF
C9343 _603_/Y _554_/A 0.59fF
C9344 _623_/X _503_/A 0.05fF
C9345 _615_/a_493_297# _593_/A 0.02fF
C9346 _387_/a_78_199# _475_/A 0.13fF
C9347 _615_/a_78_199# _593_/Y 0.38fF
C9348 _509_/Y _478_/A 0.20fF
C9349 _369_/a_76_199# _369_/a_226_297# 0.01fF
C9350 _369_/a_226_47# _369_/a_489_413# 0.02fF
C9351 _433_/Y _410_/C 0.15fF
C9352 _360_/X _361_/a_556_47# 0.02fF
C9353 _610_/A _621_/X 0.20fF
C9354 _413_/X _455_/X 0.19fF
C9355 _474_/Y _390_/B 1.21fF
C9356 _421_/a_226_47# _421_/X 0.05fF
C9357 _469_/a_664_47# _545_/Y 0.12fF
C9358 _386_/A _393_/A 0.37fF
C9359 _585_/B _381_/B 0.24fF
C9360 _385_/a_841_47# _475_/A 0.07fF
C9361 _528_/a_299_297# _557_/Y 0.01fF
C9362 VPWR _466_/X 2.76fF
C9363 _504_/X _524_/X 0.16fF
C9364 _370_/a_68_297# _370_/a_150_297# 0.02fF
C9365 _627_/A _446_/X 0.36fF
C9366 _504_/a_77_199# _471_/Y 0.15fF
C9367 _563_/a_27_297# _563_/D 0.13fF
C9368 _408_/a_68_297# VPWR 0.32fF
C9369 _433_/a_397_297# _431_/X 0.12fF
C9370 output32/a_27_47# _530_/X 0.40fF
C9371 VPWR _618_/A 3.82fF
C9372 _439_/X _510_/A 0.01fF
C9373 _342_/X _344_/a_493_297# 0.04fF
C9374 _586_/S _564_/a_27_53# 0.26fF
C9375 _359_/B VPWR 0.78fF
C9376 _353_/a_68_297# VPWR 0.35fF
C9377 _626_/Y _616_/Y 0.06fF
C9378 B[1] _368_/B 0.09fF
C9379 _540_/X _410_/C 0.01fF
C9380 _429_/a_489_413# _350_/X 0.07fF
C9381 _456_/a_76_199# VPWR 0.41fF
C9382 _559_/X _559_/a_227_47# 0.04fF
C9383 _412_/X _408_/X 0.03fF
C9384 _469_/A _571_/a_93_21# 0.15fF
C9385 _515_/Y _542_/A 0.23fF
C9386 _606_/Y _618_/A 0.21fF
C9387 _543_/Y _542_/A 1.24fF
C9388 _444_/A _390_/B 0.53fF
C9389 _510_/A _350_/C 0.20fF
C9390 _540_/a_250_297# _570_/A 0.01fF
C9391 A[5] B[4] 0.01fF
C9392 _417_/A _352_/X 0.03fF
C9393 _451_/A _514_/A 0.01fF
C9394 _447_/a_68_297# _447_/B 0.49fF
C9395 _567_/Y _469_/X 0.30fF
C9396 _423_/X _406_/Y 0.03fF
C9397 _360_/X B[1] 0.05fF
C9398 _626_/Y _550_/a_78_199# 0.13fF
C9399 _488_/a_76_199# _539_/A 0.01fF
C9400 B[0] _469_/X 0.18fF
C9401 _442_/a_27_47# _410_/C 0.22fF
C9402 _504_/a_77_199# _504_/X 0.22fF
C9403 _629_/a_68_297# _629_/a_150_297# 0.02fF
C9404 _608_/a_493_297# VPWR 0.01fF
C9405 _549_/X VPWR 2.87fF
C9406 _542_/A _521_/a_78_199# 0.01fF
C9407 _466_/X _501_/Y 0.11fF
C9408 VPWR _627_/a_27_297# 0.45fF
C9409 _584_/A _433_/Y 0.13fF
C9410 _550_/X _469_/A 0.03fF
C9411 _538_/A _539_/X 0.13fF
C9412 _533_/X _626_/Y 0.03fF
C9413 _545_/Y A[3] 0.03fF
C9414 _390_/D _520_/X 0.03fF
C9415 _487_/X _479_/a_68_297# 0.07fF
C9416 _510_/A _367_/C 0.34fF
C9417 _612_/Y _590_/A 0.14fF
C9418 _586_/S _584_/A 1.41fF
C9419 _474_/Y _471_/A 0.11fF
C9420 _419_/X _452_/A 2.84fF
C9421 _567_/B _502_/a_215_47# 0.16fF
C9422 _519_/a_29_53# _519_/A 0.57fF
C9423 _413_/X _452_/A 0.16fF
C9424 _381_/C _520_/a_76_199# 0.08fF
C9425 _542_/B _355_/A 0.44fF
C9426 _490_/X _456_/a_226_47# 0.01fF
C9427 _627_/X VPWR 1.43fF
C9428 _417_/D _519_/A 0.48fF
C9429 _378_/A _311_/a_27_47# 0.07fF
C9430 _544_/A _544_/a_381_47# 0.10fF
C9431 _485_/A _530_/X 0.08fF
C9432 _627_/A _442_/D 0.07fF
C9433 _382_/B _447_/B 0.03fF
C9434 _487_/a_78_199# _485_/D 0.00fF
C9435 _534_/a_209_297# VPWR 0.45fF
C9436 _540_/a_584_47# _472_/B 0.03fF
C9437 _386_/X _393_/A 0.21fF
C9438 _461_/a_215_47# _406_/A 0.01fF
C9439 _519_/A _332_/X 1.69fF
C9440 output17/a_27_47# _631_/Y 0.41fF
C9441 _465_/a_109_47# _427_/A 0.02fF
C9442 _419_/X _421_/X 0.22fF
C9443 _561_/A _453_/a_250_297# 0.14fF
C9444 _476_/X _472_/Y 0.78fF
C9445 _585_/B _593_/A 0.20fF
C9446 _350_/C _631_/A 0.20fF
C9447 _360_/X _383_/X 1.61fF
C9448 _318_/a_27_47# _390_/D 0.53fF
C9449 _585_/B _542_/A 1.87fF
C9450 _347_/A _541_/a_493_297# 0.13fF
C9451 _340_/A _547_/X 0.03fF
C9452 _633_/A VPWR 0.51fF
C9453 _572_/B _381_/B 0.45fF
C9454 _594_/a_27_297# _594_/X 0.23fF
C9455 B[2] _616_/A 0.38fF
C9456 _505_/a_80_21# _410_/C 0.16fF
C9457 _475_/a_68_297# _472_/B 0.07fF
C9458 _431_/a_226_47# VPWR 0.08fF
C9459 _629_/A _629_/X 0.73fF
C9460 _543_/B _417_/D 0.03fF
C9461 _313_/A _409_/a_78_199# 0.01fF
C9462 _437_/X _439_/a_76_199# 0.39fF
C9463 _410_/C _316_/a_664_47# 0.12fF
C9464 _443_/B _410_/C 0.50fF
C9465 _454_/X _449_/A 0.03fF
C9466 _588_/A _547_/X 0.20fF
C9467 _543_/B _347_/A 0.25fF
C9468 _487_/X _538_/A 0.28fF
C9469 _631_/A _367_/C 1.27fF
C9470 _406_/B _503_/A 0.58fF
C9471 input9/a_27_47# _417_/D 0.26fF
C9472 _442_/A _483_/X 0.51fF
C9473 _444_/Y _446_/a_93_21# 0.36fF
C9474 _542_/C _479_/a_68_297# 0.08fF
C9475 _343_/a_76_199# _329_/X 0.35fF
C9476 _566_/A _547_/X 0.72fF
C9477 _567_/Y _546_/X 0.24fF
C9478 _436_/X VPWR 1.01fF
C9479 _600_/a_27_297# _594_/X 0.01fF
C9480 _565_/a_209_297# _417_/D 0.14fF
C9481 _491_/X _504_/X 0.48fF
C9482 _386_/X _400_/a_80_21# 0.23fF
C9483 _469_/A _530_/X 0.03fF
C9484 _412_/X _422_/X 0.03fF
C9485 _448_/A _519_/C 0.23fF
C9486 _378_/A _584_/A 0.33fF
C9487 _318_/a_27_47# _328_/A 0.18fF
C9488 _584_/A _346_/a_161_47# 0.03fF
C9489 _422_/a_489_413# _421_/X 0.14fF
C9490 _379_/a_78_199# _419_/X 0.14fF
C9491 _487_/a_78_199# A[6] 0.05fF
C9492 _417_/D _538_/Y 0.08fF
C9493 _632_/a_292_297# _475_/A 0.06fF
C9494 _313_/a_27_47# _442_/B 0.07fF
C9495 _350_/a_109_297# _442_/B 0.01fF
C9496 _474_/Y _504_/a_77_199# 0.30fF
C9497 _576_/a_226_47# _576_/a_489_413# 0.02fF
C9498 _576_/a_76_199# _576_/a_226_297# 0.01fF
C9499 _380_/A _510_/A 0.03fF
C9500 B[2] _620_/a_226_47# 0.02fF
C9501 _596_/a_76_199# _600_/a_27_297# 0.08fF
C9502 _390_/B _430_/X 0.03fF
C9503 _503_/A _469_/a_841_47# 0.13fF
C9504 _447_/X _542_/A 0.11fF
C9505 _561_/A _514_/A 0.01fF
C9506 _591_/Y _573_/Y 0.10fF
C9507 _408_/X _631_/B 0.45fF
C9508 _328_/A _352_/a_222_93# 0.28fF
C9509 _563_/D _355_/A 0.30fF
C9510 _631_/B _320_/a_161_47# 0.01fF
C9511 A[6] _442_/A 1.22fF
C9512 _621_/a_78_199# _621_/X 0.21fF
C9513 _417_/A _542_/D 0.45fF
C9514 _430_/A _363_/B 0.02fF
C9515 _480_/A _480_/Y 1.24fF
C9516 _445_/X _443_/B 0.12fF
C9517 _424_/a_226_47# _406_/B 0.00fF
C9518 _424_/a_489_413# _406_/A 0.00fF
C9519 _466_/X _531_/C 0.01fF
C9520 _487_/X _488_/X 0.76fF
C9521 M[7] _556_/A 0.12fF
C9522 _380_/A _485_/D 0.31fF
C9523 _595_/a_227_47# _381_/B 0.01fF
C9524 _570_/X _571_/a_346_47# 0.05fF
C9525 _605_/a_80_21# _605_/a_209_47# 0.04fF
C9526 _397_/a_226_47# _397_/X 0.12fF
C9527 _436_/A _412_/X 0.28fF
C9528 _538_/A _570_/A 0.25fF
C9529 _563_/B _542_/A 2.00fF
C9530 _580_/A M[0] 0.13fF
C9531 _442_/D _316_/a_841_47# 0.03fF
C9532 _629_/A _432_/B 0.64fF
C9533 _445_/A _391_/A 0.01fF
C9534 _408_/X _411_/X 1.65fF
C9535 _569_/A _621_/X 0.08fF
C9536 B[0] _488_/a_226_47# 0.08fF
C9537 _567_/B _472_/B 0.34fF
C9538 _423_/a_493_297# VPWR 0.01fF
C9539 _572_/B _593_/A 0.02fF
C9540 _524_/a_78_199# _524_/a_292_297# 0.03fF
C9541 _474_/A VPWR 2.50fF
C9542 _516_/A _480_/A 0.01fF
C9543 _539_/a_68_297# _540_/a_93_21# 0.00fF
C9544 _493_/a_493_297# VPWR 0.01fF
C9545 _607_/a_78_199# _607_/a_215_47# 0.26fF
C9546 _480_/Y _481_/A 0.52fF
C9547 _480_/A _539_/A 0.28fF
C9548 _367_/a_27_297# _367_/a_277_297# 0.05fF
C9549 _475_/A _438_/X 0.03fF
C9550 _573_/A _573_/Y 0.74fF
C9551 M[12] VPWR 0.66fF
C9552 _417_/D _486_/X 1.62fF
C9553 _556_/Y _604_/a_303_47# 0.07fF
C9554 output24/a_27_47# _591_/A 0.28fF
C9555 _417_/A _350_/X 0.64fF
C9556 _572_/A _469_/X 0.06fF
C9557 VPWR _453_/a_250_297# 0.74fF
C9558 _380_/A _631_/A 0.09fF
C9559 _347_/A _486_/X 0.21fF
C9560 _443_/A _442_/A 0.06fF
C9561 _478_/A _466_/a_215_47# 0.11fF
C9562 _540_/a_93_21# _540_/a_250_297# 0.50fF
C9563 _513_/A _417_/D 0.89fF
C9564 _613_/X _586_/S 0.00fF
C9565 _603_/Y _579_/X 0.16fF
C9566 _390_/D _574_/X 0.16fF
C9567 _612_/Y _503_/A 0.11fF
C9568 B[2] _619_/Y 0.02fF
C9569 _469_/a_664_47# _622_/C 0.08fF
C9570 _390_/D _503_/A 0.12fF
C9571 _411_/a_68_297# _437_/a_79_199# 0.00fF
C9572 _513_/A _347_/A 0.07fF
C9573 _523_/X _492_/a_76_199# 0.01fF
C9574 _524_/a_215_47# VPWR 0.04fF
C9575 _448_/B _356_/a_215_47# 0.24fF
C9576 _627_/D _621_/X 0.37fF
C9577 _516_/A _481_/A 0.56fF
C9578 _608_/a_78_199# _469_/X 0.00fF
C9579 _542_/D _484_/a_215_47# 0.02fF
C9580 _418_/X _378_/a_558_47# 0.02fF
C9581 _481_/A _539_/A 0.47fF
C9582 _533_/X _551_/a_489_413# 0.01fF
C9583 _550_/X _551_/a_76_199# 0.23fF
C9584 _551_/X _551_/a_226_47# 0.05fF
C9585 _524_/a_78_199# _626_/Y 0.17fF
C9586 _371_/B _361_/X 0.26fF
C9587 _386_/A _505_/a_80_21# 0.16fF
C9588 _612_/Y _606_/A 0.10fF
C9589 _437_/X _402_/a_27_47# 0.18fF
C9590 _417_/D _454_/X 0.03fF
C9591 _375_/X _420_/X 0.84fF
C9592 _390_/D _606_/A 0.48fF
C9593 _384_/X B[5] 0.01fF
C9594 _386_/A _443_/B 0.30fF
C9595 _559_/X _547_/X 0.05fF
C9596 _386_/a_62_47# _570_/A 0.10fF
C9597 _575_/X _540_/X 0.01fF
C9598 _542_/D _469_/X 0.19fF
C9599 _335_/a_62_47# _335_/a_381_47# 0.08fF
C9600 _418_/B _367_/C 0.20fF
C9601 _442_/D _333_/a_27_47# 0.02fF
C9602 _336_/a_78_199# _519_/A 0.15fF
C9603 _352_/X _374_/a_215_47# 0.11fF
C9604 _455_/X _510_/A 0.11fF
C9605 _380_/A A[6] 0.05fF
C9606 _368_/B _368_/a_68_297# 0.30fF
C9607 _432_/A _432_/a_68_297# 0.50fF
C9608 _604_/X VPWR 1.16fF
C9609 _347_/A _454_/X 0.03fF
C9610 _633_/Y _489_/X 0.16fF
C9611 _542_/B _386_/a_381_47# 0.16fF
C9612 _476_/a_256_47# _469_/X 0.03fF
C9613 VPWR _394_/a_62_47# 0.52fF
C9614 _615_/a_78_199# _595_/X 0.28fF
C9615 _410_/B _433_/Y 0.03fF
C9616 _448_/A _381_/C 0.58fF
C9617 _424_/a_76_199# _433_/Y 0.08fF
C9618 _360_/X _362_/a_489_413# 0.09fF
C9619 _371_/a_68_297# _371_/B 0.41fF
C9620 _613_/X _610_/Y 0.03fF
C9621 _390_/D _549_/a_76_199# 0.07fF
C9622 _495_/a_556_47# _492_/X 0.02fF
C9623 _536_/Y _585_/B 0.46fF
C9624 _444_/A _444_/Y 1.50fF
C9625 _390_/D _390_/a_27_47# 0.46fF
C9626 _422_/X _631_/B 0.05fF
C9627 VPWR _514_/A 2.27fF
C9628 _583_/X input3/a_664_47# 0.20fF
C9629 _520_/a_226_47# _547_/a_222_93# 0.02fF
C9630 _330_/A _350_/B 0.87fF
C9631 VPWR _467_/a_397_297# 0.64fF
C9632 A[3] _622_/C 0.03fF
C9633 B[7] _449_/A 0.18fF
C9634 _587_/A _535_/Y 0.03fF
C9635 _540_/a_346_47# _410_/C 0.06fF
C9636 _347_/A _451_/A 0.11fF
C9637 _624_/a_206_369# _624_/a_489_47# 0.04fF
C9638 _623_/a_489_413# _621_/X 0.08fF
C9639 _442_/B _343_/X 0.09fF
C9640 _386_/a_62_47# _535_/A 0.02fF
C9641 _382_/A _452_/A 0.62fF
C9642 _485_/a_27_47# _484_/a_78_199# 0.00fF
C9643 input10/a_27_47# B[5] 0.07fF
C9644 M[8] _465_/a_109_297# 0.02fF
C9645 _383_/a_489_413# VPWR 0.39fF
C9646 _569_/A _568_/a_227_47# 0.18fF
C9647 _544_/A _486_/A 0.86fF
C9648 _375_/X _328_/X 0.41fF
C9649 _461_/X VPWR 5.35fF
C9650 _478_/A _469_/X 0.05fF
C9651 _546_/a_226_47# _544_/a_381_47# 0.01fF
C9652 _382_/X _420_/a_448_47# 0.14fF
C9653 _627_/C _593_/A 0.08fF
C9654 _572_/A _546_/X 0.03fF
C9655 _488_/a_76_199# _559_/X 0.02fF
C9656 _419_/X _475_/A 0.67fF
C9657 _514_/a_68_297# _515_/A 0.27fF
C9658 _457_/a_489_413# _446_/X 0.16fF
C9659 _627_/A _627_/a_27_297# 0.40fF
C9660 _360_/X _374_/a_493_297# 0.08fF
C9661 _571_/a_93_21# _570_/a_68_297# 0.00fF
C9662 _385_/a_558_47# VPWR 0.25fF
C9663 _480_/A _479_/A 0.03fF
C9664 B[7] _593_/Y 0.03fF
C9665 _390_/B _438_/X 0.83fF
C9666 _381_/C _390_/B 0.23fF
C9667 _627_/X _627_/A 0.12fF
C9668 _392_/A VPWR 2.04fF
C9669 _569_/Y _584_/A 0.08fF
C9670 _410_/B _442_/a_27_47# 0.01fF
C9671 _629_/B M[5] 1.47fF
C9672 _549_/X _548_/X 0.01fF
C9673 _439_/X _437_/X 0.09fF
C9674 _386_/X _443_/B 0.01fF
C9675 _412_/a_226_47# VPWR 0.11fF
C9676 _436_/A _631_/B 0.87fF
C9677 A[4] _427_/Y 0.07fF
C9678 _503_/a_62_47# _510_/A 0.16fF
C9679 _520_/a_226_47# _518_/X 0.25fF
C9680 _467_/a_397_297# _501_/Y 0.14fF
C9681 _420_/X _458_/a_215_47# 0.10fF
C9682 _516_/A _413_/a_68_297# 0.48fF
C9683 _623_/a_226_47# _623_/a_489_413# 0.02fF
C9684 _337_/A _332_/X 0.30fF
C9685 _371_/B _432_/X 0.11fF
C9686 _390_/D _446_/a_93_21# 0.07fF
C9687 _371_/A _430_/X 0.04fF
C9688 _407_/a_27_47# VPWR 0.03fF
C9689 _510_/A _336_/a_215_47# 0.12fF
C9690 _311_/a_27_47# _519_/A 0.24fF
C9691 _519_/X _563_/B 0.17fF
C9692 _394_/a_558_47# _394_/a_841_47# 0.07fF
C9693 _479_/A _481_/A 0.23fF
C9694 _340_/A _481_/A 0.08fF
C9695 _330_/A _384_/a_556_47# 0.02fF
C9696 _496_/a_215_47# _461_/X 0.10fF
C9697 _561_/A _512_/a_215_47# 0.20fF
C9698 _390_/D _391_/B 0.28fF
C9699 _557_/A _527_/A 0.01fF
C9700 _589_/a_76_199# A[3] 0.08fF
C9701 _360_/a_489_413# _455_/X 0.13fF
C9702 _409_/a_78_199# _445_/a_68_297# 0.02fF
C9703 _531_/B VPWR 2.65fF
C9704 _353_/X _375_/a_448_47# 0.14fF
C9705 _534_/a_80_21# _547_/X 0.10fF
C9706 _436_/A _411_/X 0.23fF
C9707 A[1] M[10] 0.16fF
C9708 _439_/X _439_/a_76_199# 0.22fF
C9709 _559_/a_323_297# _535_/Y 0.01fF
C9710 _468_/X _457_/X 0.13fF
C9711 VPWR _431_/X 1.80fF
C9712 _361_/X _361_/a_76_199# 0.29fF
C9713 _542_/C _390_/B 0.58fF
C9714 _523_/a_556_47# _522_/X 0.02fF
C9715 _417_/D _627_/B 0.01fF
C9716 _468_/X _467_/Y 0.16fF
C9717 _410_/a_197_47# VPWR 0.02fF
C9718 _411_/a_150_297# _386_/X 0.02fF
C9719 _538_/A _540_/a_93_21# 0.31fF
C9720 _516_/A _515_/Y 0.74fF
C9721 _633_/Y _588_/A 1.30fF
C9722 _390_/D _567_/a_109_297# 0.02fF
C9723 _544_/A _324_/a_62_47# 0.01fF
C9724 input12/a_62_47# input12/a_381_47# 0.08fF
C9725 _420_/X _328_/a_150_297# 0.01fF
C9726 _469_/a_558_47# VPWR 0.23fF
C9727 _440_/X VPWR 1.16fF
C9728 _432_/A _430_/a_68_297# 0.16fF
C9729 _379_/a_78_199# _382_/A 0.21fF
C9730 A[0] B[5] 0.03fF
C9731 _631_/B _350_/X 0.30fF
C9732 _335_/a_381_47# _510_/A 0.59fF
C9733 _469_/a_381_47# _469_/A 0.02fF
C9734 _564_/a_27_53# _564_/A 0.18fF
C9735 _452_/A _631_/A 0.19fF
C9736 _342_/a_68_297# _383_/X 0.14fF
C9737 _623_/a_76_199# _627_/B 0.23fF
C9738 _519_/a_29_53# _561_/A 0.20fF
C9739 VPWR _449_/A 2.42fF
C9740 _542_/C _390_/a_197_47# 0.03fF
C9741 _604_/a_80_21# _556_/A 0.12fF
C9742 _410_/B _443_/B 0.97fF
C9743 _337_/B _420_/X 0.75fF
C9744 _455_/X _443_/A 0.06fF
C9745 _417_/D _561_/A 1.33fF
C9746 _430_/A _629_/A 0.49fF
C9747 _343_/a_226_47# VPWR 0.14fF
C9748 _633_/Y _521_/a_493_297# 0.02fF
C9749 _336_/a_215_47# _631_/A 0.11fF
C9750 _518_/a_93_21# _486_/X 0.04fF
C9751 _539_/a_68_297# _483_/X 0.10fF
C9752 _442_/B _350_/B 0.16fF
C9753 _591_/Y _612_/Y 0.16fF
C9754 _520_/a_226_47# _520_/X 0.05fF
C9755 _383_/a_226_47# _383_/X 0.05fF
C9756 _347_/A _561_/A 1.24fF
C9757 _567_/B _446_/X 0.35fF
C9758 _417_/D B[7] 0.08fF
C9759 _530_/X _547_/X 6.34fF
C9760 _489_/a_489_413# _488_/X 0.16fF
C9761 _489_/a_226_297# _483_/X 0.04fF
C9762 _378_/a_381_47# VPWR 0.41fF
C9763 _585_/a_109_297# _591_/A 0.02fF
C9764 _587_/A A[3] 0.10fF
C9765 _442_/a_303_47# _478_/A 0.03fF
C9766 _584_/a_68_297# _584_/A 0.32fF
C9767 _612_/A A[3] 0.24fF
C9768 _330_/A _371_/B 0.03fF
C9769 _614_/a_489_413# output24/a_27_47# 0.03fF
C9770 _567_/B _532_/a_206_369# 0.05fF
C9771 B[1] _313_/A 0.03fF
C9772 _530_/X _570_/a_68_297# 0.07fF
C9773 VPWR _593_/Y 5.12fF
C9774 _440_/a_76_199# _440_/a_489_413# 0.12fF
C9775 _416_/a_78_199# _324_/a_381_47# 0.05fF
C9776 _507_/a_109_297# _507_/Y 0.03fF
C9777 _463_/a_226_47# VPWR 0.05fF
C9778 _322_/A _355_/A 0.07fF
C9779 _538_/Y _410_/C 0.25fF
C9780 _584_/A _564_/A 0.01fF
C9781 _392_/Y VPWR 1.46fF
C9782 _568_/a_77_199# _543_/Y 0.02fF
C9783 _385_/a_664_47# _393_/A 0.10fF
C9784 input3/a_841_47# VPWR 0.31fF
C9785 _568_/a_227_297# _567_/B 0.09fF
C9786 _432_/A _629_/a_68_297# 0.20fF
C9787 _585_/B _539_/A 0.84fF
C9788 VPWR _554_/B 1.85fF
C9789 _539_/a_68_297# A[6] 0.15fF
C9790 _455_/X _418_/B 0.02fF
C9791 _625_/Y A[3] 0.15fF
C9792 _537_/a_227_297# _472_/B 0.03fF
C9793 _416_/a_78_199# _378_/A 0.13fF
C9794 _527_/Y _527_/A 0.80fF
C9795 _503_/A _631_/Y 0.08fF
C9796 _570_/B _469_/X 1.38fF
C9797 _551_/X M[0] 0.45fF
C9798 _436_/A _349_/a_493_297# 0.08fF
C9799 _611_/X _621_/a_215_47# 0.03fF
C9800 _506_/Y _442_/A 1.11fF
C9801 _384_/a_226_297# _384_/a_76_199# 0.01fF
C9802 _466_/a_292_297# _431_/X 0.01fF
C9803 output31/a_27_47# _464_/A 0.02fF
C9804 _466_/a_78_199# _432_/X 0.30fF
C9805 VPWR _575_/a_292_297# 0.01fF
C9806 _378_/A M[9] 0.07fF
C9807 _516_/A _386_/a_841_47# 0.05fF
C9808 _457_/a_76_199# _457_/X 0.22fF
C9809 _512_/a_215_47# VPWR 0.06fF
C9810 _328_/B _419_/X 0.03fF
C9811 M[5] _399_/a_78_199# 0.04fF
C9812 _543_/A _442_/D 0.03fF
C9813 _610_/A _590_/B 1.33fF
C9814 _387_/a_215_47# _391_/A 0.01fF
C9815 _569_/Y _613_/X 0.10fF
C9816 _515_/Y _340_/A 0.04fF
C9817 _503_/a_381_47# _503_/A 0.02fF
C9818 _576_/a_226_297# _574_/X 0.01fF
C9819 _444_/A _390_/D 0.45fF
C9820 _475_/X _472_/B 0.99fF
C9821 _445_/A _563_/D 0.45fF
C9822 _572_/a_68_297# _585_/B 0.08fF
C9823 _368_/B _633_/Y 0.01fF
C9824 _410_/C _486_/X 0.69fF
C9825 B[0] _479_/B 0.22fF
C9826 _567_/B _498_/Y 0.50fF
C9827 _342_/X _343_/a_226_47# 0.01fF
C9828 _437_/a_79_199# _437_/a_448_47# 0.13fF
C9829 _439_/a_226_47# _438_/X 0.53fF
C9830 _633_/Y _559_/X 0.03fF
C9831 output27/a_27_47# _373_/a_113_297# 0.02fF
C9832 M[2] VPWR 1.67fF
C9833 _440_/a_226_47# _439_/X 0.52fF
C9834 _543_/Y _588_/A 0.11fF
C9835 _630_/a_76_199# VPWR 0.46fF
C9836 _513_/A _410_/C 0.11fF
C9837 _360_/X _481_/A 0.53fF
C9838 _498_/A VPWR 2.05fF
C9839 _464_/A _626_/Y 0.20fF
C9840 _566_/A _515_/Y 0.02fF
C9841 _566_/A _543_/Y 1.56fF
C9842 _360_/X _633_/Y 0.12fF
C9843 _452_/A _418_/B 0.22fF
C9844 _568_/a_77_199# _585_/B 0.03fF
C9845 _519_/a_29_53# VPWR 0.53fF
C9846 _510_/A _510_/X 0.23fF
C9847 _607_/X _616_/Y 0.23fF
C9848 _381_/B _469_/X 0.59fF
C9849 _586_/a_76_199# _586_/a_218_374# 0.03fF
C9850 _417_/D VPWR 6.12fF
C9851 _520_/a_76_199# A[6] 0.05fF
C9852 _409_/a_215_47# _481_/A 0.22fF
C9853 _607_/a_215_47# _606_/A 0.07fF
C9854 _543_/B _386_/A 0.24fF
C9855 _347_/A VPWR 6.61fF
C9856 _531_/B _531_/C 0.73fF
C9857 _454_/X _410_/C 1.30fF
C9858 VPWR _332_/X 1.63fF
C9859 _538_/A _485_/D 0.09fF
C9860 M[2] _314_/X 0.07fF
C9861 _371_/B _442_/B 0.03fF
C9862 _417_/A _542_/A 0.22fF
C9863 _570_/B _546_/X 0.10fF
C9864 _362_/a_76_199# _361_/X 0.22fF
C9865 _464_/A _406_/Y 0.18fF
C9866 _547_/a_222_93# _486_/B 0.21fF
C9867 _623_/a_76_199# VPWR 0.49fF
C9868 _565_/a_209_297# _386_/A 0.22fF
C9869 _318_/a_27_47# _326_/A 0.02fF
C9870 _429_/a_489_413# _363_/B 0.11fF
C9871 _433_/Y _535_/Y 0.05fF
C9872 _351_/X _361_/a_226_47# 0.01fF
C9873 _584_/A _486_/X 0.20fF
C9874 _386_/a_381_47# _520_/X 0.08fF
C9875 _547_/X _514_/B 0.19fF
C9876 input9/a_27_47# _521_/X 0.16fF
C9877 _384_/X _384_/a_76_199# 0.22fF
C9878 _530_/a_489_413# VPWR 0.36fF
C9879 _503_/a_381_47# _471_/Y 0.01fF
C9880 _469_/a_62_47# _469_/X 0.49fF
C9881 _586_/a_505_21# _622_/C 0.24fF
C9882 _510_/A _475_/A 2.68fF
C9883 _533_/X _539_/A 0.01fF
C9884 _513_/A _584_/A 0.07fF
C9885 _538_/A _483_/X 0.02fF
C9886 _459_/a_226_47# _459_/a_489_413# 0.02fF
C9887 _506_/A _505_/a_80_21# 0.20fF
C9888 _624_/a_206_369# _624_/X 0.04fF
C9889 _585_/B _588_/A 0.32fF
C9890 _536_/a_109_297# VPWR 0.01fF
C9891 _444_/A _389_/a_27_47# 0.10fF
C9892 _411_/B _412_/X 0.00fF
C9893 _374_/a_78_199# _361_/X 0.36fF
C9894 _406_/Y _631_/B 0.04fF
C9895 _540_/X _535_/Y 0.12fF
C9896 _533_/X _489_/X 0.27fF
C9897 _566_/A _585_/B 0.07fF
C9898 _542_/a_27_47# _515_/A 0.01fF
C9899 M[2] _342_/X 0.03fF
C9900 _591_/A _622_/C 1.23fF
C9901 _626_/Y _523_/a_76_199# 0.08fF
C9902 _572_/a_68_297# _572_/B 0.59fF
C9903 _518_/X _486_/B 0.02fF
C9904 _584_/A _454_/X 0.03fF
C9905 _525_/a_489_413# _524_/X 0.14fF
C9906 _353_/X _519_/A 0.53fF
C9907 _542_/A _484_/a_215_47# 0.02fF
C9908 _328_/B _335_/a_62_47# 0.00fF
C9909 _433_/Y _432_/X 0.55fF
C9910 _444_/Y _542_/C 0.20fF
C9911 _516_/A _322_/a_27_47# 0.02fF
C9912 _381_/B _546_/X 0.16fF
C9913 _569_/A _570_/X 0.28fF
C9914 _542_/A _469_/X 0.05fF
C9915 _386_/A _486_/X 0.17fF
C9916 _557_/Y _583_/a_76_199# 0.01fF
C9917 _524_/a_215_47# _523_/X 0.08fF
C9918 _400_/a_209_297# _392_/Y 0.23fF
C9919 _400_/a_80_21# _330_/A 0.18fF
C9920 _583_/a_226_47# _582_/Y 0.59fF
C9921 _583_/a_76_199# _602_/A 0.37fF
C9922 _483_/X _488_/X 2.83fF
C9923 _451_/A _584_/A 0.26fF
C9924 _469_/a_664_47# _433_/Y 0.10fF
C9925 _554_/X _491_/X 0.00fF
C9926 B[1] _408_/B 0.12fF
C9927 _487_/a_292_297# _519_/C 0.02fF
C9928 _331_/a_27_47# _350_/B 0.47fF
C9929 _487_/a_215_47# _449_/A 0.11fF
C9930 input3/a_381_47# input3/a_558_47# 0.32fF
C9931 _469_/a_664_47# _586_/S 0.02fF
C9932 _469_/a_558_47# _627_/A 0.19fF
C9933 _563_/A _449_/A 0.31fF
C9934 _386_/a_558_47# _386_/A 0.08fF
C9935 _432_/B input14/a_27_47# 0.01fF
C9936 _454_/a_76_199# _454_/a_489_413# 0.12fF
C9937 _475_/A _631_/A 0.64fF
C9938 _580_/A _551_/X 0.35fF
C9939 _329_/a_226_47# _442_/B 0.14fF
C9940 _513_/A _386_/A 0.53fF
C9941 _555_/a_215_297# _556_/A 0.15fF
C9942 _448_/B _481_/A 0.14fF
C9943 input9/a_27_47# _550_/a_215_47# 0.03fF
C9944 _551_/a_226_47# _551_/a_489_413# 0.02fF
C9945 _551_/a_76_199# _551_/a_226_297# 0.01fF
C9946 _455_/X _506_/Y 0.47fF
C9947 _616_/A _599_/Y 0.03fF
C9948 _598_/a_68_297# _616_/A 0.24fF
C9949 _512_/a_78_199# _542_/A 0.04fF
C9950 _535_/Y _537_/a_539_297# 0.02fF
C9951 _520_/X _522_/X 0.62fF
C9952 _509_/Y _539_/A 0.05fF
C9953 _506_/Y _509_/A 0.03fF
C9954 _633_/a_74_47# _631_/A 0.00fF
C9955 _558_/a_77_199# _558_/a_227_47# 0.24fF
C9956 _545_/Y _503_/A 0.41fF
C9957 _603_/Y _604_/X 0.00fF
C9958 B[6] _401_/A 0.24fF
C9959 _398_/a_226_47# _374_/X 0.25fF
C9960 _633_/Y _530_/X 0.03fF
C9961 _386_/A _454_/X 0.03fF
C9962 M[1] _442_/D 0.06fF
C9963 B[7] _624_/a_76_199# 0.20fF
C9964 _537_/a_77_199# _410_/C 0.00fF
C9965 _564_/a_219_297# _622_/X 0.00fF
C9966 _564_/a_27_53# _627_/B 0.05fF
C9967 A[6] _488_/X 0.08fF
C9968 _522_/X _522_/a_489_413# 0.00fF
C9969 _359_/a_68_297# _454_/X 0.11fF
C9970 _561_/A _311_/a_27_47# 0.10fF
C9971 _502_/a_78_199# _502_/a_215_47# 0.26fF
C9972 _510_/A _473_/a_77_199# 0.38fF
C9973 _526_/a_76_199# _504_/X 0.47fF
C9974 _588_/A _572_/B 0.27fF
C9975 _390_/D _539_/X 0.16fF
C9976 _500_/a_78_199# _427_/A 0.01fF
C9977 _443_/A _443_/a_68_297# 0.38fF
C9978 _422_/a_76_199# VPWR 0.50fF
C9979 _408_/B _383_/X 0.03fF
C9980 _510_/A _390_/B 0.65fF
C9981 _375_/X B[1] 0.28fF
C9982 _423_/a_292_297# _396_/X 0.08fF
C9983 _512_/a_78_199# _512_/a_292_297# 0.03fF
C9984 M[1] _588_/Y 0.07fF
C9985 _381_/C _381_/a_303_47# 0.06fF
C9986 _498_/A _531_/C 0.22fF
C9987 input13/a_27_47# VPWR 0.52fF
C9988 _393_/A _442_/B 0.17fF
C9989 _566_/A _572_/B 0.18fF
C9990 _477_/a_78_199# VPWR 0.60fF
C9991 _525_/a_76_199# VPWR 0.45fF
C9992 _386_/X _486_/X 0.21fF
C9993 _454_/a_489_413# _447_/X 0.07fF
C9994 _454_/a_226_47# _453_/X 0.56fF
C9995 _583_/a_76_199# _606_/A 0.08fF
C9996 _336_/a_78_199# VPWR 0.63fF
C9997 _441_/a_78_199# _355_/A 0.37fF
C9998 _444_/A _631_/Y 0.23fF
C9999 _386_/a_558_47# _386_/X 0.25fF
C10000 _595_/X VPWR 4.35fF
C10001 A[4] _427_/A 0.01fF
C10002 A[3] _540_/X 0.27fF
C10003 _590_/A _622_/C 0.65fF
C10004 VPWR _518_/a_93_21# 0.39fF
C10005 _584_/A _627_/B 1.76fF
C10006 _583_/X _442_/D 5.78fF
C10007 _627_/D _590_/B 0.03fF
C10008 _494_/a_76_199# _494_/a_226_47# 0.49fF
C10009 output20/a_27_47# M[12] 0.41fF
C10010 _587_/A _591_/A 0.27fF
C10011 _382_/a_68_297# _383_/a_76_199# 0.03fF
C10012 _396_/X input14/a_27_47# 0.00fF
C10013 _583_/X _579_/X 0.36fF
C10014 _485_/A _517_/X 0.01fF
C10015 _612_/A _591_/A 0.10fF
C10016 _366_/a_76_199# _366_/a_226_47# 0.49fF
C10017 _442_/D _622_/X 0.17fF
C10018 _378_/a_558_47# _324_/a_381_47# 0.01fF
C10019 B[0] _542_/D 0.03fF
C10020 _487_/X _486_/A 0.25fF
C10021 _436_/A _408_/X 1.37fF
C10022 _596_/a_226_47# VPWR 0.10fF
C10023 _461_/a_78_199# _424_/X 0.28fF
C10024 _371_/B _397_/X 0.03fF
C10025 _491_/X _525_/a_489_413# 0.10fF
C10026 _490_/X _525_/a_226_47# 0.01fF
C10027 _380_/A _350_/C 0.04fF
C10028 _614_/a_76_199# M[1] 0.01fF
C10029 _544_/A _565_/a_80_21# 0.10fF
C10030 _328_/B _510_/A 0.91fF
C10031 _330_/A _351_/a_219_297# 0.06fF
C10032 _396_/a_93_21# _392_/A 0.31fF
C10033 _588_/a_109_297# VPWR 0.01fF
C10034 _375_/X _383_/X 2.22fF
C10035 VPWR _547_/a_79_199# 0.65fF
C10036 _534_/a_80_21# _515_/Y 0.18fF
C10037 _386_/X _454_/X 0.03fF
C10038 _544_/A _545_/Y 0.21fF
C10039 _519_/A M[9] 0.83fF
C10040 _575_/a_78_199# _547_/X 0.13fF
C10041 _360_/X _359_/X 0.57fF
C10042 output25/a_27_47# M[2] 0.44fF
C10043 _619_/a_27_47# _607_/a_215_47# 0.06fF
C10044 _510_/X _472_/Y 0.17fF
C10045 _510_/A _471_/A 0.05fF
C10046 _601_/Y _607_/a_78_199# 0.01fF
C10047 _487_/X _390_/D 1.57fF
C10048 _561_/A _584_/A 0.13fF
C10049 _587_/A _624_/a_206_369# 0.01fF
C10050 _336_/a_78_199# _314_/X 0.03fF
C10051 _597_/a_493_297# _575_/X 0.08fF
C10052 _597_/a_78_199# _598_/B 0.25fF
C10053 _597_/a_215_47# _576_/X 0.05fF
C10054 _458_/X _457_/X 2.51fF
C10055 _411_/B _411_/X 0.80fF
C10056 _625_/Y _591_/A 0.11fF
C10057 _595_/a_227_47# _588_/A 0.09fF
C10058 _623_/X _621_/X 1.01fF
C10059 _417_/D _563_/A 0.39fF
C10060 _519_/X _484_/a_215_47# 0.02fF
C10061 VPWR _462_/a_226_297# 0.00fF
C10062 B[7] _584_/A 0.53fF
C10063 _445_/X _446_/a_584_47# 0.01fF
C10064 input5/a_62_47# _478_/A 0.31fF
C10065 _381_/C _486_/A 0.13fF
C10066 _524_/a_78_199# _489_/X 0.01fF
C10067 _497_/B _464_/A 0.11fF
C10068 _347_/A _563_/A 0.06fF
C10069 VPWR _624_/a_76_199# 0.53fF
C10070 _417_/D _627_/A 0.05fF
C10071 _380_/A _442_/A 0.35fF
C10072 _577_/a_226_47# VPWR 0.12fF
C10073 _554_/X _555_/a_215_297# 0.06fF
C10074 _390_/D _381_/C 0.61fF
C10075 _569_/Y _571_/a_250_297# 0.04fF
C10076 _625_/Y _624_/a_206_369# 0.01fF
C10077 _544_/A _447_/B 1.12fF
C10078 _513_/A _410_/B 0.01fF
C10079 _627_/C _588_/A 0.12fF
C10080 _404_/a_381_47# _404_/a_841_47# 0.03fF
C10081 _404_/a_558_47# _404_/a_664_47# 0.60fF
C10082 _625_/a_27_297# _625_/a_277_47# 0.04fF
C10083 _543_/Y _530_/X 0.06fF
C10084 _581_/a_27_93# _602_/A 0.35fF
C10085 _515_/Y _530_/X 0.29fF
C10086 _461_/a_215_47# _390_/B 0.02fF
C10087 _494_/a_76_199# _493_/X 0.24fF
C10088 _563_/D _393_/A 0.39fF
C10089 _567_/B _436_/X 0.34fF
C10090 _602_/Y _530_/X 0.25fF
C10091 _366_/a_76_199# _337_/X 0.25fF
C10092 _311_/a_27_47# VPWR 0.66fF
C10093 _459_/X _458_/X 1.29fF
C10094 _328_/B _631_/A 1.25fF
C10095 _391_/a_68_297# _391_/a_150_297# 0.02fF
C10096 M[2] _368_/A 0.19fF
C10097 input10/a_27_47# _398_/X 0.00fF
C10098 VPWR _410_/C 7.29fF
C10099 _623_/X _623_/a_226_47# 0.05fF
C10100 _455_/X _359_/A 0.20fF
C10101 _458_/X _503_/A 0.03fF
C10102 _390_/D _570_/A 0.05fF
C10103 _329_/a_76_199# _338_/X 0.02fF
C10104 _410_/B _454_/X 1.41fF
C10105 _456_/a_226_47# _454_/X 0.25fF
C10106 _442_/A _316_/a_381_47# 0.02fF
C10107 _550_/a_292_297# _550_/a_78_199# 0.03fF
C10108 _442_/A _508_/a_227_297# 0.04fF
C10109 _410_/B _334_/a_27_47# 0.36fF
C10110 _390_/D _316_/a_62_47# 0.18fF
C10111 _564_/a_27_53# VPWR 0.13fF
C10112 _616_/Y _616_/B 0.45fF
C10113 _589_/a_489_413# _588_/Y 0.14fF
C10114 _542_/C _390_/D 0.45fF
C10115 _436_/X _468_/a_78_199# 0.38fF
C10116 _443_/A _390_/B 0.03fF
C10117 _578_/a_78_199# _578_/a_215_47# 0.26fF
C10118 M[12] input12/a_841_47# 0.05fF
C10119 _544_/A _486_/a_68_297# 0.29fF
C10120 _504_/a_77_199# _510_/A 0.36fF
C10121 _598_/B _601_/A 0.35fF
C10122 _442_/B _332_/a_150_297# 0.01fF
C10123 VPWR _507_/a_109_297# 0.01fF
C10124 _587_/A _520_/X 0.04fF
C10125 _633_/Y _385_/a_381_47# 0.08fF
C10126 _332_/X _368_/A 0.52fF
C10127 _603_/Y _554_/B 0.75fF
C10128 _631_/B _337_/X 0.42fF
C10129 _426_/A _466_/X 0.04fF
C10130 _587_/A _590_/A 0.34fF
C10131 _572_/B _571_/a_93_21# 0.13fF
C10132 _568_/a_323_297# VPWR 0.02fF
C10133 _353_/X _337_/A 0.12fF
C10134 _590_/A _612_/A 0.27fF
C10135 _390_/D _535_/A 0.03fF
C10136 _453_/X _542_/D 0.03fF
C10137 _506_/A _507_/Y 0.10fF
C10138 _396_/a_93_21# _392_/Y 0.34fF
C10139 _519_/C _628_/Y 0.01fF
C10140 _585_/B _530_/X 0.49fF
C10141 _445_/X VPWR 0.74fF
C10142 _442_/a_27_47# _442_/B 0.29fF
C10143 B[7] _454_/a_556_47# 0.02fF
C10144 _542_/a_27_47# _542_/B 0.27fF
C10145 M[10] _558_/X 0.51fF
C10146 _583_/X _611_/X 0.01fF
C10147 _406_/A _421_/X 0.12fF
C10148 _420_/a_544_297# VPWR 0.01fF
C10149 _584_/A VPWR 9.34fF
C10150 _607_/X B[2] 0.59fF
C10151 _455_/X _442_/A 5.39fF
C10152 _429_/a_226_47# _398_/a_226_47# 0.01fF
C10153 _602_/Y _557_/B 0.20fF
C10154 _533_/a_77_199# _539_/A 0.30fF
C10155 _399_/a_292_297# _398_/X 0.08fF
C10156 _420_/a_79_199# VPWR 0.73fF
C10157 _415_/a_27_47# _561_/A 0.31fF
C10158 _359_/A _452_/A 0.01fF
C10159 _625_/Y _590_/A 0.32fF
C10160 _608_/a_78_199# _572_/A 0.06fF
C10161 _374_/a_78_199# _442_/B 0.13fF
C10162 _496_/a_78_199# _460_/X 0.01fF
C10163 _397_/X _399_/a_493_297# 0.08fF
C10164 _503_/A _622_/C 1.07fF
C10165 _516_/A _417_/A 0.40fF
C10166 VPWR _522_/a_226_47# 0.06fF
C10167 _410_/B _337_/A 0.02fF
C10168 _594_/a_27_297# _593_/Y 0.32fF
C10169 _513_/A _485_/a_27_47# 0.13fF
C10170 _313_/A _481_/A 0.01fF
C10171 _348_/a_27_47# _408_/B 0.31fF
C10172 _550_/X _550_/a_78_199# 0.20fF
C10173 _322_/A _441_/a_215_47# 0.16fF
C10174 _318_/a_27_47# _326_/a_27_47# 0.01fF
C10175 _572_/A _542_/D 0.03fF
C10176 _417_/a_109_47# VPWR 0.00fF
C10177 _313_/A _633_/Y 0.58fF
C10178 _492_/a_226_47# VPWR 0.11fF
C10179 _533_/X _550_/X 0.26fF
C10180 _418_/B _418_/A 0.46fF
C10181 _452_/X _519_/C 1.35fF
C10182 _510_/X _506_/Y 0.51fF
C10183 _499_/a_384_47# _497_/A 0.13fF
C10184 _419_/X _632_/a_215_47# 0.02fF
C10185 _609_/a_209_297# _622_/C 0.24fF
C10186 input5/a_664_47# VPWR 0.33fF
C10187 _626_/a_481_47# _612_/A 0.01fF
C10188 _389_/a_27_47# _316_/a_62_47# 0.01fF
C10189 _523_/a_76_199# _523_/a_226_47# 0.49fF
C10190 _473_/a_77_199# _472_/Y 0.42fF
C10191 _583_/X _618_/A 1.18fF
C10192 _626_/Y _599_/Y 0.99fF
C10193 _600_/a_27_297# _593_/Y 0.02fF
C10194 _542_/C _389_/a_27_47# 0.22fF
C10195 _620_/a_76_199# _620_/a_489_413# 0.12fF
C10196 _608_/a_78_199# _542_/D 0.00fF
C10197 _563_/D _586_/S 0.00fF
C10198 _485_/a_303_47# A[6] 0.03fF
C10199 _330_/A _351_/A 1.53fF
C10200 _549_/a_76_199# _549_/a_226_297# 0.01fF
C10201 _549_/a_226_47# _549_/a_489_413# 0.02fF
C10202 _419_/X _328_/A 0.03fF
C10203 _618_/Y _606_/A 0.15fF
C10204 _613_/X B[7] 0.53fF
C10205 _447_/X _530_/X 0.00fF
C10206 _556_/Y _602_/Y 0.91fF
C10207 _532_/a_76_199# _527_/Y 0.30fF
C10208 B[7] _575_/X 0.34fF
C10209 _595_/a_227_47# _571_/a_93_21# 0.06fF
C10210 _626_/a_397_297# VPWR 0.52fF
C10211 _352_/a_79_199# VPWR 0.55fF
C10212 _567_/Y _570_/B 0.74fF
C10213 _544_/A _486_/B 0.33fF
C10214 _488_/a_226_47# _488_/a_489_413# 0.02fF
C10215 _488_/a_76_199# _488_/a_226_297# 0.01fF
C10216 _548_/a_489_413# _547_/X 0.29fF
C10217 _548_/a_226_47# _546_/X 0.33fF
C10218 _538_/A _559_/a_77_199# 0.05fF
C10219 _452_/A _367_/C 0.05fF
C10220 _527_/B _528_/a_299_297# 0.25fF
C10221 _562_/a_78_199# _562_/a_215_47# 0.26fF
C10222 _316_/a_62_47# _316_/a_558_47# 0.03fF
C10223 B[0] _626_/Y 0.02fF
C10224 _508_/a_77_199# _508_/a_323_297# 0.05fF
C10225 _626_/a_481_47# _625_/Y 0.07fF
C10226 _386_/A VPWR 4.20fF
C10227 _442_/B _443_/B 0.18fF
C10228 _543_/B _515_/A 0.12fF
C10229 _543_/A _514_/A 0.54fF
C10230 _543_/Y _514_/B 0.11fF
C10231 _542_/B _443_/B 0.14fF
C10232 _557_/B _558_/a_227_297# 0.07fF
C10233 M[2] _370_/A 0.09fF
C10234 _628_/a_28_47# _627_/X 0.21fF
C10235 _613_/X _589_/a_226_47# 0.02fF
C10236 _515_/Y _514_/B 0.04fF
C10237 _359_/a_68_297# VPWR 0.27fF
C10238 _358_/a_27_47# _485_/A 0.64fF
C10239 _469_/A _521_/a_215_47# 0.20fF
C10240 _444_/A _443_/a_150_297# 0.01fF
C10241 _336_/a_215_47# _367_/C 0.12fF
C10242 _436_/A _350_/X 0.37fF
C10243 _569_/Y A[3] 2.57fF
C10244 _387_/a_78_199# _313_/a_27_47# 0.00fF
C10245 VPWR _398_/a_489_413# 0.32fF
C10246 _384_/X _631_/A 0.34fF
C10247 _431_/a_226_47# _426_/A 0.09fF
C10248 VPWR _521_/X 1.30fF
C10249 _455_/X _380_/A 0.83fF
C10250 _614_/a_226_47# VPWR 0.08fF
C10251 _608_/a_215_47# _627_/B 0.10fF
C10252 _440_/X _460_/a_226_47# 0.31fF
C10253 _468_/X _438_/X 0.01fF
C10254 _419_/X _421_/a_226_297# 0.05fF
C10255 _539_/A _469_/X 0.38fF
C10256 _586_/a_505_21# _433_/Y 0.12fF
C10257 _342_/a_150_297# _420_/X 0.01fF
C10258 _482_/a_68_297# _482_/a_150_297# 0.02fF
C10259 _513_/A _506_/A 0.03fF
C10260 _627_/A _595_/X 0.06fF
C10261 _352_/a_79_199# _314_/X 0.01fF
C10262 _614_/a_226_297# _623_/X 0.02fF
C10263 _539_/a_68_297# _442_/A 0.07fF
C10264 _605_/a_303_47# _557_/Y 0.05fF
C10265 VPWR _483_/a_93_21# 0.41fF
C10266 _337_/a_68_297# _338_/X 0.16fF
C10267 _582_/Y VPWR 1.26fF
C10268 _586_/S _586_/a_505_21# 0.38fF
C10269 _454_/a_556_47# VPWR 0.00fF
C10270 _432_/a_68_297# _432_/a_150_297# 0.02fF
C10271 _626_/Y _492_/X 0.46fF
C10272 _472_/Y _471_/A 0.08fF
C10273 _545_/Y _546_/a_226_47# 0.70fF
C10274 _360_/a_76_199# VPWR 0.34fF
C10275 _419_/a_76_199# _419_/X 0.22fF
C10276 _610_/A _621_/a_78_199# 0.25fF
C10277 _533_/X _530_/X 0.52fF
C10278 _557_/A output30/a_27_47# 0.19fF
C10279 _413_/X _419_/a_76_199# 0.40fF
C10280 _620_/a_226_47# _619_/Y 0.55fF
C10281 _381_/C _628_/Y 0.40fF
C10282 _447_/a_68_297# _519_/A 0.20fF
C10283 _375_/a_222_93# _455_/X 0.13fF
C10284 _461_/a_292_297# VPWR 0.01fF
C10285 _567_/Y _381_/B 0.08fF
C10286 _487_/X _452_/X 0.01fF
C10287 _415_/a_27_47# VPWR 0.49fF
C10288 B[0] _381_/B 0.10fF
C10289 _416_/a_215_47# _418_/B 0.12fF
C10290 _563_/D _346_/a_161_47# 0.13fF
C10291 _538_/Y _535_/Y 0.77fF
C10292 _392_/A _420_/X 0.37fF
C10293 _495_/a_76_199# _497_/A 0.22fF
C10294 _569_/A _610_/A 0.03fF
C10295 _487_/X _481_/a_27_47# 0.07fF
C10296 _387_/a_78_199# _326_/A 0.00fF
C10297 _426_/A _373_/a_199_47# 0.01fF
C10298 _557_/B _558_/X 0.28fF
C10299 _567_/B _531_/B 0.03fF
C10300 _359_/B _485_/A 0.00fF
C10301 _587_/A _503_/A 2.93fF
C10302 _338_/a_222_93# _332_/X 0.03fF
C10303 _595_/a_227_297# _566_/Y 0.01fF
C10304 _342_/X _352_/a_79_199# 0.17fF
C10305 _595_/a_77_199# _570_/X 0.28fF
C10306 _386_/X VPWR 4.64fF
C10307 _612_/A _503_/A 0.02fF
C10308 _591_/Y _624_/X 0.04fF
C10309 _427_/Y _464_/Y 0.36fF
C10310 _381_/C _452_/X 0.31fF
C10311 _432_/A _629_/B 1.24fF
C10312 _343_/X B[5] 0.18fF
C10313 _613_/X VPWR 3.03fF
C10314 _426_/a_68_297# VPWR 0.34fF
C10315 _382_/B _519_/A 0.03fF
C10316 _515_/A _486_/X 0.16fF
C10317 VPWR _550_/a_215_47# 0.07fF
C10318 _563_/B _453_/a_93_21# 0.01fF
C10319 _543_/B _469_/a_664_47# 0.02fF
C10320 _543_/A _469_/a_558_47# 0.01fF
C10321 _575_/X VPWR 3.82fF
C10322 _440_/X _567_/B 0.57fF
C10323 _631_/B _328_/a_68_297# 0.08fF
C10324 _563_/A _410_/C 0.13fF
C10325 _611_/a_109_297# _592_/a_113_297# 0.01fF
C10326 _386_/a_558_47# _515_/A 0.14fF
C10327 input7/a_27_47# _489_/a_76_199# 0.02fF
C10328 _631_/Y _316_/a_62_47# 0.10fF
C10329 _428_/a_299_297# _427_/Y 0.05fF
C10330 _338_/a_448_47# _337_/X 0.22fF
C10331 _542_/C _631_/Y 0.80fF
C10332 _615_/a_292_297# _593_/Y 0.02fF
C10333 _544_/a_558_47# _503_/A 0.03fF
C10334 _475_/A _402_/a_27_47# 0.01fF
C10335 _446_/a_93_21# _446_/a_346_47# 0.05fF
C10336 _610_/A _627_/D 0.74fF
C10337 _387_/a_292_297# _475_/A 0.02fF
C10338 _548_/a_76_199# _548_/a_226_47# 0.49fF
C10339 _353_/X VPWR 2.27fF
C10340 _335_/a_62_47# _328_/A 0.15fF
C10341 _610_/Y _591_/A 0.44fF
C10342 _599_/A _576_/X 0.00fF
C10343 _416_/a_78_199# _561_/A 0.47fF
C10344 _556_/Y _558_/X 0.01fF
C10345 VPWR _609_/a_80_21# 0.40fF
C10346 _535_/Y _486_/X 0.00fF
C10347 _631_/Y _552_/a_226_47# 0.01fF
C10348 _350_/a_27_297# _350_/C 0.55fF
C10349 _380_/a_27_47# _442_/A 0.21fF
C10350 _591_/Y _622_/C 0.19fF
C10351 _598_/a_68_297# _593_/A 0.01fF
C10352 _525_/X _524_/X 1.11fF
C10353 _561_/A M[9] 0.07fF
C10354 _481_/a_27_47# _570_/A 0.01fF
C10355 _433_/a_397_297# _432_/X 0.12fF
C10356 _342_/X _344_/a_215_47# 0.06fF
C10357 _586_/S _564_/a_301_297# 0.01fF
C10358 _601_/Y _606_/A 0.79fF
C10359 M[8] _390_/B 0.41fF
C10360 _497_/A _468_/X 0.52fF
C10361 _626_/Y _616_/A 0.40fF
C10362 _474_/A _476_/a_93_21# 0.34fF
C10363 _503_/A _559_/a_323_297# 0.05fF
C10364 _410_/B VPWR 4.96fF
C10365 _429_/a_226_297# _350_/X 0.04fF
C10366 _525_/a_76_199# _523_/X 0.41fF
C10367 _424_/a_76_199# VPWR 0.58fF
C10368 _475_/X _436_/X 0.01fF
C10369 A[3] _507_/Y 0.48fF
C10370 _587_/A _471_/Y 1.39fF
C10371 _476_/X _390_/B 0.01fF
C10372 _588_/A _469_/X 0.73fF
C10373 _570_/B _572_/A 0.18fF
C10374 B[0] _542_/A 0.70fF
C10375 _408_/B _633_/Y 0.03fF
C10376 _544_/A _587_/A 0.12fF
C10377 _419_/X _631_/Y 0.03fF
C10378 _447_/a_150_297# _447_/B 0.02fF
C10379 _388_/a_27_47# _390_/B 0.02fF
C10380 _566_/A _469_/X 0.47fF
C10381 _340_/A _512_/a_78_199# 0.42fF
C10382 _573_/A _622_/C 0.03fF
C10383 _422_/X _406_/Y 0.25fF
C10384 _563_/A _584_/A 1.41fF
C10385 _424_/X _461_/X 0.01fF
C10386 _583_/X M[12] 0.28fF
C10387 _442_/a_109_47# _410_/C 0.04fF
C10388 _445_/X _470_/a_80_21# 0.01fF
C10389 _382_/a_68_297# _382_/a_150_297# 0.02fF
C10390 _580_/B VPWR 0.93fF
C10391 _520_/X _433_/Y 0.13fF
C10392 _488_/a_226_47# _539_/A 0.02fF
C10393 _358_/a_27_47# _383_/X 0.23fF
C10394 M[10] _501_/a_397_297# 0.03fF
C10395 _513_/A _381_/a_27_47# 0.31fF
C10396 _608_/a_215_47# VPWR 0.11fF
C10397 _375_/X _396_/X 0.05fF
C10398 _519_/C _447_/B 0.17fF
C10399 _382_/X _419_/X 0.51fF
C10400 _590_/A _433_/Y 0.13fF
C10401 _487_/X _479_/a_150_297# 0.01fF
C10402 VPWR _590_/a_68_297# 0.33fF
C10403 _633_/Y _472_/B 1.59fF
C10404 _376_/X VPWR 1.81fF
C10405 _586_/S _590_/A 0.29fF
C10406 _627_/A _584_/A 0.70fF
C10407 _568_/a_77_199# _546_/X 0.13fF
C10408 _392_/Y _420_/X 0.30fF
C10409 _452_/a_68_297# _452_/a_150_297# 0.02fF
C10410 _411_/B _408_/X 0.04fF
C10411 _519_/a_111_297# _519_/A 0.03fF
C10412 _442_/D M[6] 0.23fF
C10413 _455_/X _452_/A 0.03fF
C10414 _542_/C _355_/A 0.43fF
C10415 _544_/A _544_/a_558_47# 0.14fF
C10416 _635_/Y B[5] 0.62fF
C10417 _482_/a_68_297# _539_/A 0.30fF
C10418 _538_/Y A[3] 0.14fF
C10419 _482_/X _483_/a_584_47# 0.01fF
C10420 B[2] _559_/X 0.62fF
C10421 _633_/A _367_/a_27_297# 0.00fF
C10422 _520_/X _540_/X 0.58fF
C10423 _440_/a_76_199# _458_/X 0.07fF
C10424 _587_/A _566_/Y 0.37fF
C10425 _375_/X _481_/A 0.01fF
C10426 _461_/a_215_47# _406_/B 0.01fF
C10427 _424_/X _407_/a_27_47# 0.01fF
C10428 _380_/a_27_47# _380_/A 0.39fF
C10429 _461_/a_78_199# _407_/Y 0.37fF
C10430 _485_/D _486_/A 0.60fF
C10431 _375_/X _633_/Y 0.03fF
C10432 _475_/A _350_/C 0.83fF
C10433 _474_/A _475_/X 0.02fF
C10434 _395_/X VPWR 0.65fF
C10435 _360_/X _417_/A 0.03fF
C10436 _442_/D _547_/X 0.03fF
C10437 _318_/a_109_47# _390_/D 0.04fF
C10438 _441_/a_78_199# _441_/a_215_47# 0.26fF
C10439 _390_/D _485_/D 1.46fF
C10440 _347_/A _541_/a_215_47# 0.10fF
C10441 _594_/a_27_297# _595_/X 0.18fF
C10442 _594_/a_109_297# _594_/X 0.03fF
C10443 B[2] _616_/B 0.03fF
C10444 _519_/A _442_/B 0.88fF
C10445 _505_/a_209_297# _410_/C 0.29fF
C10446 _416_/a_78_199# VPWR 0.58fF
C10447 _437_/X _439_/a_226_47# 0.22fF
C10448 _458_/a_78_199# _458_/a_215_47# 0.26fF
C10449 _475_/A _367_/C 0.34fF
C10450 _431_/a_489_413# VPWR 0.39fF
C10451 _567_/B _417_/D 0.05fF
C10452 _359_/B _383_/X 0.35fF
C10453 _510_/A _328_/A 1.06fF
C10454 _363_/A _630_/a_76_199# 0.02fF
C10455 _513_/A _382_/B 0.05fF
C10456 _386_/A _470_/a_80_21# 0.18fF
C10457 _588_/A _546_/X 0.39fF
C10458 _445_/A _387_/a_78_199# 0.28fF
C10459 A[3] _486_/X 0.19fF
C10460 _543_/A _347_/A 0.01fF
C10461 _485_/a_27_47# VPWR 0.73fF
C10462 _444_/Y _446_/a_250_297# 0.03fF
C10463 _390_/D _483_/X 0.03fF
C10464 _557_/A _530_/X 0.03fF
C10465 _591_/Y _587_/A 0.64fF
C10466 VPWR M[9] 1.30fF
C10467 _343_/a_226_47# _329_/X 0.25fF
C10468 _600_/a_27_297# _595_/X 0.01fF
C10469 _566_/A _546_/X 1.27fF
C10470 _605_/a_80_21# _604_/a_209_297# 0.01fF
C10471 _476_/X _524_/X 0.10fF
C10472 _386_/X _400_/a_209_297# 0.22fF
C10473 _406_/A _390_/B 0.03fF
C10474 _426_/A _431_/X 0.30fF
C10475 _520_/X _537_/a_539_297# 0.04fF
C10476 _432_/A M[5] 0.32fF
C10477 VPWR M[14] 0.55fF
C10478 _587_/a_27_47# _587_/A 0.38fF
C10479 _382_/B _454_/X 0.40fF
C10480 _382_/A _419_/a_76_199# 0.01fF
C10481 _439_/a_76_199# _439_/a_226_47# 0.49fF
C10482 _621_/X _628_/Y 0.50fF
C10483 _629_/B _371_/A 0.38fF
C10484 _613_/X _613_/a_77_199# 0.22fF
C10485 _596_/a_226_47# _600_/a_27_297# 0.01fF
C10486 _350_/a_205_297# _442_/B 0.01fF
C10487 _632_/a_493_297# _475_/A 0.08fF
C10488 _420_/X _332_/X 0.03fF
C10489 B[2] _620_/a_489_413# 0.07fF
C10490 _543_/B _542_/B 0.05fF
C10491 _406_/Y _478_/A 0.13fF
C10492 A[6] _486_/A 0.35fF
C10493 _453_/X _542_/A 0.03fF
C10494 _390_/B _428_/X 0.23fF
C10495 _627_/D _621_/a_78_199# 0.12fF
C10496 B[1] _633_/A 0.04fF
C10497 _328_/A _352_/a_544_297# 0.06fF
C10498 _632_/a_215_47# _631_/A 0.23fF
C10499 _537_/a_77_199# _535_/Y 0.38fF
C10500 _591_/Y _625_/Y 0.08fF
C10501 _621_/a_493_297# _591_/A 0.01fF
C10502 _626_/a_481_47# _610_/Y 0.01fF
C10503 _390_/D A[6] 0.05fF
C10504 _587_/A _573_/A 0.73fF
C10505 _370_/B B[5] 0.39fF
C10506 _474_/Y _587_/A 0.78fF
C10507 _616_/A _593_/A 0.03fF
C10508 _439_/X _390_/B 0.43fF
C10509 _381_/C _447_/B 0.57fF
C10510 _482_/a_68_297# _479_/A 0.01fF
C10511 _318_/a_197_47# _380_/A 0.03fF
C10512 _347_/A _411_/A 0.00fF
C10513 _623_/X _590_/B 0.18fF
C10514 _455_/X _380_/a_27_47# 0.10fF
C10515 _328_/A _631_/A 0.03fF
C10516 _605_/a_80_21# _605_/a_303_47# 0.04fF
C10517 _569_/A _627_/D 0.11fF
C10518 _478_/A _381_/B 0.18fF
C10519 input3/a_664_47# _616_/Y 0.00fF
C10520 input3/a_558_47# _616_/A 0.01fF
C10521 input3/a_62_47# _618_/A 0.00fF
C10522 _462_/a_76_199# _462_/a_226_47# 0.49fF
C10523 _572_/A _593_/A 0.13fF
C10524 _623_/a_226_47# _628_/Y 0.01fF
C10525 _368_/B _366_/a_76_199# 0.00fF
C10526 _423_/a_215_47# VPWR 0.04fF
C10527 B[0] _562_/a_493_297# 0.04fF
C10528 _386_/X _470_/a_80_21# 0.01fF
C10529 _390_/B _350_/C 0.33fF
C10530 _493_/a_215_47# VPWR 0.07fF
C10531 _571_/a_93_21# _469_/X 0.21fF
C10532 M[2] _374_/X 0.01fF
C10533 _506_/A VPWR 3.70fF
C10534 _544_/a_62_47# _544_/a_381_47# 0.08fF
C10535 _567_/Y _536_/Y 0.04fF
C10536 _380_/A _475_/A 1.23fF
C10537 _557_/A _557_/B 1.35fF
C10538 _322_/A _346_/a_161_47# 0.01fF
C10539 _533_/a_227_47# _539_/A 0.02fF
C10540 _431_/a_76_199# _466_/a_215_47# 0.01fF
C10541 _362_/a_556_47# _352_/X 0.02fF
C10542 _371_/B B[5] 1.13fF
C10543 _503_/A _433_/Y 1.94fF
C10544 _393_/A _391_/B 0.14fF
C10545 _540_/a_93_21# _540_/a_256_47# 0.03fF
C10546 _417_/A _448_/B 1.03fF
C10547 _379_/a_78_199# _452_/A 0.38fF
C10548 _411_/a_68_297# _437_/a_222_93# 0.02fF
C10549 _410_/a_27_47# _478_/A 0.01fF
C10550 _527_/Y _530_/X 0.29fF
C10551 _586_/S _503_/A 0.50fF
C10552 M[2] _329_/X 0.42fF
C10553 _619_/a_27_47# _601_/Y 0.18fF
C10554 B[2] _530_/X 0.59fF
C10555 _375_/a_79_199# _376_/a_68_297# 0.00fF
C10556 _411_/a_68_297# _510_/A 0.20fF
C10557 _554_/X _583_/a_76_199# 0.01fF
C10558 _417_/A _530_/X 0.16fF
C10559 _533_/X _551_/a_226_297# 0.02fF
C10560 _386_/A _505_/a_209_297# 0.11fF
C10561 _542_/A _542_/D 1.43fF
C10562 _549_/X _551_/a_76_199# 0.34fF
C10563 _550_/X _551_/a_226_47# 0.66fF
C10564 _588_/A _548_/a_76_199# 0.00fF
C10565 M[10] _531_/A 0.01fF
C10566 _368_/B _631_/B 0.00fF
C10567 _627_/A _609_/a_80_21# 0.20fF
C10568 _386_/a_381_47# _570_/A 0.08fF
C10569 _464_/A _465_/X 0.06fF
C10570 _559_/X _546_/X 0.04fF
C10571 _542_/B _486_/X 0.03fF
C10572 _574_/X _540_/X 0.46fF
C10573 _503_/A _540_/X 0.18fF
C10574 _575_/X _548_/X 0.01fF
C10575 _335_/a_62_47# _335_/a_558_47# 0.03fF
C10576 _448_/a_68_297# _519_/C 0.01fF
C10577 _418_/A _367_/C 0.28fF
C10578 _336_/a_292_297# _519_/A 0.02fF
C10579 _557_/a_109_297# _557_/Y 0.02fF
C10580 _328_/B _350_/C 0.35fF
C10581 _404_/a_62_47# _609_/a_80_21# 0.04fF
C10582 _455_/X _510_/X 0.26fF
C10583 _557_/A _556_/Y 0.12fF
C10584 _410_/B _563_/A 0.03fF
C10585 VPWR _361_/X 0.94fF
C10586 _503_/a_841_47# _446_/X 0.07fF
C10587 VPWR _571_/a_250_297# 0.74fF
C10588 _513_/A _542_/B 0.68fF
C10589 _343_/a_76_199# _369_/a_226_47# 0.01fF
C10590 _476_/a_346_47# _469_/X 0.07fF
C10591 _585_/B _472_/B 0.74fF
C10592 VPWR _394_/a_381_47# 0.31fF
C10593 _510_/X _509_/A 0.07fF
C10594 _615_/a_292_297# _595_/X 0.08fF
C10595 _410_/B _470_/a_80_21# 0.27fF
C10596 _511_/a_93_21# _509_/A 0.39fF
C10597 _360_/X _631_/B 0.03fF
C10598 _476_/X _491_/X 2.79fF
C10599 _424_/a_226_47# _433_/Y 0.14fF
C10600 _390_/D _549_/a_226_47# 0.07fF
C10601 _400_/a_80_21# _391_/B 0.57fF
C10602 _496_/a_78_199# _496_/a_292_297# 0.03fF
C10603 _633_/Y _446_/X 1.08fF
C10604 _347_/A _409_/a_78_199# 0.14fF
C10605 _425_/a_489_413# _461_/X 0.01fF
C10606 _413_/X _447_/B 0.03fF
C10607 _478_/a_27_47# _410_/C 0.03fF
C10608 _630_/a_76_199# _426_/A 0.07fF
C10609 _328_/B _367_/C 0.17fF
C10610 VPWR _515_/A 2.34fF
C10611 _382_/A _382_/X 0.05fF
C10612 _553_/a_78_199# _554_/B 0.24fF
C10613 _559_/a_77_199# _559_/a_227_297# 0.13fF
C10614 _542_/B _454_/X 0.03fF
C10615 _540_/a_584_47# _410_/C 0.02fF
C10616 _458_/X _438_/X 0.29fF
C10617 _623_/a_226_297# _621_/X 0.03fF
C10618 _487_/X _486_/B 0.19fF
C10619 _571_/a_93_21# _546_/X 0.04fF
C10620 _494_/a_76_199# _495_/a_76_199# 0.01fF
C10621 _626_/Y _467_/a_109_47# 0.12fF
C10622 _546_/a_76_199# VPWR 0.49fF
C10623 _371_/a_68_297# VPWR 0.28fF
C10624 _510_/A _631_/Y 0.03fF
C10625 _471_/Y _433_/Y 0.48fF
C10626 _610_/A _601_/A 0.02fF
C10627 _549_/a_76_199# _540_/X 0.32fF
C10628 _608_/a_215_47# _627_/A 0.11fF
C10629 _546_/a_226_47# _544_/a_558_47# 0.05fF
C10630 _546_/a_76_199# _544_/a_664_47# 0.01fF
C10631 _488_/a_226_47# _559_/X 0.01fF
C10632 _490_/a_215_47# _446_/X 0.03fF
C10633 _530_/X _531_/A 0.06fF
C10634 _544_/A _433_/Y 0.04fF
C10635 _457_/a_226_297# _446_/X 0.01fF
C10636 VPWR _535_/Y 1.84fF
C10637 _423_/a_493_297# _383_/X 0.08fF
C10638 _360_/X _374_/a_215_47# 0.10fF
C10639 _626_/Y _406_/Y 0.23fF
C10640 _480_/Y _479_/B 0.06fF
C10641 _385_/a_664_47# VPWR 0.40fF
C10642 _530_/X _469_/X 0.03fF
C10643 _375_/X _359_/X 0.36fF
C10644 _569_/Y _590_/A 0.07fF
C10645 _380_/A _390_/B 0.66fF
C10646 _351_/A _384_/a_489_413# 0.09fF
C10647 _418_/B _324_/a_62_47# 0.24fF
C10648 _412_/a_489_413# VPWR 0.39fF
C10649 B[7] A[3] 0.17fF
C10650 _581_/B _555_/a_215_297# 0.00fF
C10651 _439_/X _504_/a_77_199# 0.00fF
C10652 _520_/a_489_413# _518_/X 0.07fF
C10653 VPWR input1/a_27_47# 0.51fF
C10654 _442_/D _481_/A 0.03fF
C10655 _516_/A _413_/a_150_297# 0.01fF
C10656 _390_/D _446_/a_250_297# 0.11fF
C10657 _428_/a_81_21# _426_/B 0.02fF
C10658 _570_/B _381_/B 0.35fF
C10659 _371_/B _430_/X 0.16fF
C10660 _373_/Y _432_/X 0.59fF
C10661 _394_/a_664_47# _394_/a_841_47# 0.29fF
C10662 _479_/B _539_/A 0.03fF
C10663 _516_/A _479_/B 0.20fF
C10664 _464_/Y _427_/A 1.37fF
C10665 _633_/Y _442_/D 0.02fF
C10666 _563_/D _486_/X 0.23fF
C10667 _452_/X _485_/D 0.01fF
C10668 B[7] M[15] 0.16fF
C10669 _607_/X _599_/Y 0.41fF
C10670 B[0] _480_/Y 0.05fF
C10671 _381_/a_27_47# VPWR 0.74fF
C10672 _562_/a_215_47# _563_/B 0.02fF
C10673 _416_/a_215_47# _367_/C 0.04fF
C10674 _526_/a_76_199# _527_/B 0.22fF
C10675 _534_/a_209_297# _547_/X 0.14fF
C10676 _439_/X _439_/a_226_47# 0.05fF
C10677 VPWR _432_/X 2.62fF
C10678 _513_/A _563_/D 0.07fF
C10679 _598_/a_68_297# _598_/A 0.32fF
C10680 _544_/A _542_/a_27_47# 0.39fF
C10681 M[2] _369_/a_76_199# 0.09fF
C10682 _631_/Y _631_/A 0.14fF
C10683 _393_/A B[5] 0.02fF
C10684 _599_/Y _598_/A 0.09fF
C10685 _567_/Y _435_/a_27_47# 0.01fF
C10686 _538_/A _540_/a_250_297# 0.05fF
C10687 _391_/A VPWR 0.99fF
C10688 _410_/a_303_47# VPWR 0.01fF
C10689 _396_/a_93_21# _386_/X 0.23fF
C10690 _633_/Y _588_/Y 0.48fF
C10691 input12/a_62_47# input12/a_558_47# 0.03fF
C10692 B[1] _392_/A 0.11fF
C10693 _381_/C _448_/a_68_297# 0.07fF
C10694 _452_/A _475_/A 0.00fF
C10695 _528_/a_81_21# _528_/a_299_297# 0.21fF
C10696 _469_/a_664_47# VPWR 0.35fF
C10697 _516_/A B[0] 0.39fF
C10698 B[0] _539_/A 0.11fF
C10699 _432_/A _430_/a_150_297# 0.02fF
C10700 _447_/a_68_297# VPWR 0.29fF
C10701 _335_/a_558_47# _510_/A 0.11fF
C10702 A[6] _628_/Y 0.03fF
C10703 _515_/Y _517_/X 0.63fF
C10704 _563_/D _454_/X 0.03fF
C10705 _342_/a_150_297# _383_/X 0.02fF
C10706 _473_/a_227_47# _472_/B 0.13fF
C10707 _567_/a_109_297# _540_/X 0.01fF
C10708 _519_/X _542_/D 0.16fF
C10709 _481_/a_27_47# _483_/X 0.01fF
C10710 _350_/B _384_/a_76_199# 0.09fF
C10711 _623_/a_76_199# _622_/X 0.27fF
C10712 _544_/A _378_/A 1.12fF
C10713 _604_/a_209_297# _556_/A 0.13fF
C10714 _542_/C _390_/a_303_47# 0.06fF
C10715 _633_/Y _521_/a_215_47# 0.02fF
C10716 _343_/a_489_413# VPWR 0.42fF
C10717 _587_/A _539_/X 0.01fF
C10718 _518_/a_250_297# _486_/X 0.21fF
C10719 _451_/a_27_47# _628_/Y 0.07fF
C10720 _530_/X _546_/X 1.31fF
C10721 _387_/a_78_199# _387_/a_215_47# 0.26fF
C10722 _611_/a_27_297# _591_/A 0.35fF
C10723 _511_/X _509_/A 0.71fF
C10724 _630_/X _350_/X 0.11fF
C10725 _476_/a_250_297# _472_/B 0.26fF
C10726 _382_/B VPWR 1.84fF
C10727 _584_/a_68_297# _590_/A 0.27fF
C10728 _612_/Y _590_/B 0.18fF
C10729 _530_/X _570_/a_150_297# 0.01fF
C10730 _440_/a_226_47# _440_/a_489_413# 0.02fF
C10731 _440_/a_76_199# _440_/a_226_297# 0.01fF
C10732 _463_/a_489_413# VPWR 0.42fF
C10733 _459_/a_226_297# _457_/X 0.04fF
C10734 _626_/Y _593_/A 0.03fF
C10735 _533_/X _554_/A 0.31fF
C10736 VPWR A[3] 3.17fF
C10737 _330_/A VPWR 4.41fF
C10738 _343_/a_489_413# _314_/X 0.01fF
C10739 _419_/X _418_/X 0.05fF
C10740 _399_/a_78_199# _399_/a_292_297# 0.03fF
C10741 _568_/a_77_199# _567_/Y 0.39fF
C10742 _568_/a_323_297# _567_/B 0.09fF
C10743 _474_/Y _433_/Y 0.11fF
C10744 _432_/A _629_/a_150_297# 0.01fF
C10745 _413_/X _418_/X 2.02fF
C10746 _599_/A _593_/Y 0.01fF
C10747 _539_/a_150_297# A[6] 0.02fF
C10748 _419_/X _395_/a_68_297# 0.01fF
C10749 _410_/B _333_/a_27_47# 0.24fF
C10750 _537_/a_323_297# _472_/B 0.11fF
C10751 _520_/X _507_/Y 0.21fF
C10752 _436_/A _349_/a_215_47# 0.22fF
C10753 _479_/B _479_/A 0.42fF
C10754 M[2] _634_/Y 0.32fF
C10755 _613_/X _621_/a_215_47# 0.21fF
C10756 _407_/Y _461_/X 0.12fF
C10757 _443_/B _446_/a_93_21# 0.15fF
C10758 _358_/a_27_47# _481_/A 0.05fF
C10759 _466_/a_493_297# _431_/X 0.01fF
C10760 VPWR M[15] 1.08fF
C10761 _466_/a_78_199# _430_/X 0.15fF
C10762 _419_/X _350_/B 0.06fF
C10763 _591_/Y _610_/Y 0.28fF
C10764 VPWR _575_/a_493_297# 0.01fF
C10765 _509_/Y _472_/B 0.15fF
C10766 _338_/X _343_/X 0.53fF
C10767 _487_/X _587_/A 0.07fF
C10768 input9/a_27_47# _520_/X 0.01fF
C10769 _632_/a_78_199# VPWR 0.57fF
C10770 _412_/a_76_199# _412_/X 0.22fF
C10771 _516_/a_27_47# _386_/X 0.17fF
C10772 _533_/a_227_297# _503_/A 0.03fF
C10773 _598_/a_68_297# _598_/a_150_297# 0.02fF
C10774 _457_/a_226_47# _457_/X 0.05fF
C10775 _350_/X _363_/B 0.94fF
C10776 _562_/a_215_47# _627_/C 0.20fF
C10777 _515_/Y _442_/D 0.41fF
C10778 _543_/Y _442_/D 0.18fF
C10779 _518_/X _486_/X 0.17fF
C10780 _455_/a_79_199# _416_/a_78_199# 0.02fF
C10781 _444_/Y _442_/A 0.28fF
C10782 _569_/Y _503_/A 0.54fF
C10783 _455_/X _471_/A 0.01fF
C10784 _467_/Y _500_/a_215_47# 0.02fF
C10785 input5/a_62_47# input5/a_381_47# 0.08fF
C10786 _513_/A _518_/X 0.80fF
C10787 _356_/a_78_199# _359_/A 0.21fF
C10788 _390_/D _559_/a_77_199# 0.19fF
C10789 B[0] _479_/A 0.33fF
C10790 _503_/a_62_47# _473_/a_77_199# 0.01fF
C10791 B[0] _340_/A 0.12fF
C10792 _611_/X _633_/Y 0.34fF
C10793 _600_/a_285_47# _616_/B 0.04fF
C10794 _587_/A _438_/X 0.46fF
C10795 _457_/X _460_/a_76_199# 0.08fF
C10796 _497_/a_68_297# _497_/a_150_297# 0.02fF
C10797 _407_/a_27_47# _407_/Y 0.29fF
C10798 _406_/A _406_/B 0.87fF
C10799 _538_/Y _520_/X 0.12fF
C10800 _437_/a_222_93# _437_/a_448_47# 0.03fF
C10801 _439_/a_489_413# _438_/X 0.14fF
C10802 _420_/a_79_199# _420_/X 0.37fF
C10803 _440_/a_489_413# _439_/X 0.14fF
C10804 _630_/a_226_47# VPWR 0.09fF
C10805 _623_/X _610_/A 0.15fF
C10806 _396_/a_93_21# _395_/X 0.22fF
C10807 _567_/Y _588_/A 0.43fF
C10808 _381_/B _542_/A 0.39fF
C10809 _445_/X _411_/A 0.01fF
C10810 _367_/a_27_297# _332_/X 0.01fF
C10811 _454_/X _518_/X 0.51fF
C10812 _567_/Y _566_/A 0.41fF
C10813 _519_/a_111_297# VPWR 0.00fF
C10814 _452_/A _418_/A 0.84fF
C10815 _510_/X _511_/a_93_21# 0.25fF
C10816 _566_/A B[0] 0.03fF
C10817 _607_/X _616_/A 0.21fF
C10818 _520_/a_226_47# A[6] 0.06fF
C10819 _380_/A _361_/a_226_47# 0.00fF
C10820 _548_/a_76_199# _530_/X 0.17fF
C10821 _417_/D _469_/A 0.11fF
C10822 _421_/a_76_199# VPWR 0.48fF
C10823 A[7] _376_/X 0.08fF
C10824 _587_/A _570_/A 0.18fF
C10825 _359_/B _481_/A 0.35fF
C10826 _351_/a_219_297# B[5] 0.08fF
C10827 _443_/A _355_/A 0.01fF
C10828 _327_/a_78_199# _335_/a_62_47# 0.02fF
C10829 _440_/X _459_/a_76_199# 0.06fF
C10830 _497_/B _626_/Y 1.28fF
C10831 _351_/X _371_/B 0.55fF
C10832 _611_/a_27_297# _590_/A 0.01fF
C10833 _616_/A _598_/A 0.27fF
C10834 _444_/A _442_/a_27_47# 0.02fF
C10835 M[0] _530_/X 0.11fF
C10836 _563_/D _561_/A 0.59fF
C10837 _487_/X _559_/a_323_297# 0.03fF
C10838 _459_/X _460_/a_76_199# 0.25fF
C10839 _513_/a_27_47# _543_/Y 0.14fF
C10840 _362_/a_226_47# _361_/X 0.53fF
C10841 _464_/A _462_/X 0.01fF
C10842 _569_/A _595_/a_77_199# 0.06fF
C10843 _346_/A _340_/a_27_47# 0.00fF
C10844 _520_/X _486_/X 2.71fF
C10845 _456_/a_76_199# _633_/Y 0.08fF
C10846 _392_/Y _383_/X 0.00fF
C10847 _429_/a_226_297# _363_/B 0.01fF
C10848 output26/a_27_47# A[0] 0.09fF
C10849 _410_/a_27_47# _411_/B 0.19fF
C10850 _628_/a_382_297# _621_/X 0.02fF
C10851 _521_/a_78_199# _521_/a_215_47# 0.26fF
C10852 _386_/a_558_47# _520_/X 0.08fF
C10853 _580_/A _559_/X 0.03fF
C10854 _342_/a_68_297# _631_/B 0.39fF
C10855 _503_/a_62_47# _471_/A 0.10fF
C10856 _503_/a_381_47# _472_/Y 0.01fF
C10857 _328_/B _336_/a_215_47# 0.01fF
C10858 _530_/a_226_297# VPWR 0.00fF
C10859 _384_/X _384_/a_226_47# 0.05fF
C10860 _442_/B VPWR 7.87fF
C10861 _542_/B VPWR 3.54fF
C10862 _555_/a_27_413# _555_/a_215_297# 0.43fF
C10863 _577_/a_76_199# _533_/X 0.02fF
C10864 _485_/D _447_/B 0.43fF
C10865 _500_/a_215_47# _427_/A 0.16fF
C10866 _469_/a_381_47# _469_/X 0.69fF
C10867 _355_/a_161_47# _584_/A 0.03fF
C10868 _497_/B _406_/Y 0.20fF
C10869 M[4] _373_/Y 0.06fF
C10870 _506_/A _505_/a_209_297# 0.04fF
C10871 _445_/A _335_/a_62_47# 0.58fF
C10872 _587_/A _535_/A 0.41fF
C10873 VPWR _552_/a_76_199# 0.46fF
C10874 _456_/a_76_199# _490_/a_215_47# 0.01fF
C10875 _506_/A _508_/a_227_47# 0.05fF
C10876 _506_/Y _508_/a_323_297# 0.06fF
C10877 _386_/A _411_/A 0.52fF
C10878 _542_/C _514_/a_68_297# 0.00fF
C10879 _602_/Y _558_/a_227_47# 0.01fF
C10880 M[4] VPWR 0.52fF
C10881 _621_/X _622_/C 0.06fF
C10882 _626_/Y _523_/a_226_47# 0.11fF
C10883 _572_/a_68_297# _572_/A 0.33fF
C10884 _363_/A _344_/a_215_47# 0.01fF
C10885 input7/a_27_47# _521_/a_78_199# 0.02fF
C10886 _488_/a_556_47# _469_/A 0.05fF
C10887 _525_/a_226_297# _524_/X 0.01fF
C10888 _352_/a_79_199# _328_/X 0.27fF
C10889 _628_/a_382_297# _623_/a_226_47# 0.01fF
C10890 _314_/X _442_/B 1.18fF
C10891 _563_/A _391_/A 0.21fF
C10892 _444_/A _443_/B 1.38fF
C10893 _445_/X _409_/a_78_199# 0.01fF
C10894 _380_/a_27_47# _390_/B 0.02fF
C10895 _412_/a_76_199# _631_/B 0.07fF
C10896 _465_/a_27_297# _464_/Y 0.14fF
C10897 input4/a_27_47# _542_/A 0.07fF
C10898 _423_/a_215_47# _396_/a_93_21# 0.09fF
C10899 _524_/a_78_199# _554_/A 0.00fF
C10900 _569_/Y _566_/Y 0.49fF
C10901 _416_/a_215_47# _452_/A 0.07fF
C10902 _417_/a_27_47# _447_/X 0.03fF
C10903 _485_/D _486_/a_68_297# 0.19fF
C10904 _503_/A _507_/Y 0.17fF
C10905 _400_/a_209_297# _330_/A 0.09fF
C10906 _615_/a_215_47# _616_/B 0.01fF
C10907 _634_/a_27_413# VPWR 0.28fF
C10908 _583_/a_489_413# _582_/Y 0.14fF
C10909 _583_/a_226_47# _602_/A 0.34fF
C10910 _543_/B _503_/A 0.01fF
C10911 _628_/a_300_47# _564_/a_219_297# 0.03fF
C10912 _487_/a_493_297# _519_/C 0.02fF
C10913 input3/a_381_47# input3/a_664_47# 0.09fF
C10914 _567_/Y _559_/X 0.48fF
C10915 _386_/a_664_47# _386_/A 0.31fF
C10916 _454_/a_76_199# _454_/a_226_297# 0.01fF
C10917 _454_/a_226_47# _454_/a_489_413# 0.02fF
C10918 _633_/A _633_/Y 0.13fF
C10919 _513_/A _322_/A 0.15fF
C10920 _469_/a_664_47# _627_/A 0.28fF
C10921 _318_/a_27_47# _334_/a_27_47# 0.05fF
C10922 _555_/a_298_297# _556_/A 0.04fF
C10923 B[7] _591_/A 0.93fF
C10924 _478_/A _539_/A 0.43fF
C10925 _386_/X _420_/X 0.80fF
C10926 _412_/a_76_199# _411_/X 0.25fF
C10927 _633_/a_74_47# _475_/A 0.01fF
C10928 _344_/a_78_199# _344_/a_292_297# 0.03fF
C10929 _493_/X _460_/X 0.00fF
C10930 _598_/a_150_297# _616_/A 0.02fF
C10931 _616_/B _599_/Y 0.48fF
C10932 _535_/Y _537_/a_227_47# 0.07fF
C10933 _452_/a_68_297# _453_/a_93_21# 0.02fF
C10934 _544_/A _379_/a_493_297# 0.04fF
C10935 _342_/X _442_/B 0.29fF
C10936 _487_/a_78_199# _487_/a_292_297# 0.03fF
C10937 _586_/a_76_199# _622_/C 0.74fF
C10938 _588_/A _616_/A 0.02fF
C10939 _398_/a_489_413# _374_/X 0.07fF
C10940 _390_/D _350_/C 0.06fF
C10941 B[7] _624_/a_206_369# 0.07fF
C10942 _322_/A _454_/X 0.23fF
C10943 _630_/X output28/a_27_47# 0.46fF
C10944 _563_/D VPWR 4.37fF
C10945 _510_/X _511_/X 0.01fF
C10946 _386_/X _411_/A 0.39fF
C10947 _564_/a_27_53# _622_/X 0.01fF
C10948 _564_/a_301_297# _627_/B 0.01fF
C10949 _519_/X _381_/B 0.33fF
C10950 _550_/a_78_199# _522_/a_76_199# 0.04fF
C10951 _327_/a_78_199# _510_/A 0.07fF
C10952 _544_/A _519_/A 0.03fF
C10953 _522_/X _522_/a_226_297# 0.01fF
C10954 _444_/Y _455_/X 0.34fF
C10955 _359_/a_150_297# _454_/X 0.01fF
C10956 _538_/Y _503_/A 0.54fF
C10957 output17/a_27_47# VPWR 0.62fF
C10958 _511_/a_93_21# _511_/X 0.13fF
C10959 _433_/Y _539_/X 0.04fF
C10960 _353_/X _420_/X 0.24fF
C10961 _429_/a_76_199# _397_/X 0.08fF
C10962 _626_/a_109_47# _616_/A 0.09fF
C10963 _533_/X _522_/a_76_199# 0.07fF
C10964 _510_/A _473_/a_227_297# 0.04fF
C10965 _526_/a_76_199# _525_/X 0.22fF
C10966 _526_/a_226_47# _504_/X 0.22fF
C10967 _463_/a_76_199# _464_/A 0.24fF
C10968 _417_/A _408_/B 0.35fF
C10969 input12/a_62_47# _618_/Y 0.01fF
C10970 _442_/D _620_/a_76_199# 0.03fF
C10971 _628_/a_28_47# _584_/A 0.12fF
C10972 _588_/A _572_/A 1.14fF
C10973 _485_/A _547_/a_79_199# 0.12fF
C10974 _427_/Y VPWR 1.91fF
C10975 _422_/a_226_47# VPWR 0.09fF
C10976 _610_/A _469_/a_841_47# 0.03fF
C10977 _350_/C _332_/a_68_297# 0.17fF
C10978 _506_/Y _631_/Y 0.18fF
C10979 _536_/Y _381_/B 0.05fF
C10980 _525_/a_226_47# VPWR 0.06fF
C10981 _477_/a_292_297# VPWR 0.01fF
C10982 _627_/A A[3] 0.09fF
C10983 _384_/X _397_/a_76_199# 0.37fF
C10984 _627_/C _564_/a_219_297# 0.11fF
C10985 _390_/D _442_/A 0.12fF
C10986 _375_/X _329_/a_556_47# 0.02fF
C10987 A[2] _390_/D 0.06fF
C10988 _540_/X _539_/X 0.45fF
C10989 _390_/B _443_/a_68_297# 0.01fF
C10990 _454_/a_226_297# _447_/X 0.02fF
C10991 _454_/a_489_413# _453_/X 0.14fF
C10992 _616_/a_109_297# VPWR 0.01fF
C10993 _576_/a_76_199# VPWR 0.54fF
C10994 _583_/a_226_47# _606_/A 0.14fF
C10995 _336_/a_292_297# VPWR 0.01fF
C10996 _445_/A _510_/A 0.83fF
C10997 _583_/X _584_/A 0.01fF
C10998 _632_/a_215_47# _367_/C 0.03fF
C10999 _344_/a_215_47# _329_/X 0.11fF
C11000 _569_/A _623_/X 0.03fF
C11001 _587_/A _540_/a_93_21# 0.01fF
C11002 _386_/a_664_47# _386_/X 0.15fF
C11003 _485_/D _486_/B 0.31fF
C11004 _544_/A _543_/B 2.16fF
C11005 _351_/A B[5] 0.11fF
C11006 _586_/a_505_21# VPWR 0.34fF
C11007 _584_/A _622_/X 0.27fF
C11008 _520_/X _537_/a_77_199# 0.13fF
C11009 _505_/a_80_21# _482_/X 0.29fF
C11010 VPWR _518_/a_250_297# 0.70fF
C11011 _428_/a_81_21# _428_/X 0.24fF
C11012 _410_/B _511_/a_346_47# 0.02fF
C11013 _590_/A _627_/B 0.24fF
C11014 _580_/A _530_/X 1.19fF
C11015 _503_/A _486_/X 0.06fF
C11016 _494_/a_76_199# _494_/a_489_413# 0.12fF
C11017 _382_/a_68_297# _383_/a_226_47# 0.01fF
C11018 _474_/A _633_/Y 0.03fF
C11019 _360_/X _352_/X 3.76fF
C11020 _558_/a_227_47# _558_/X 0.04fF
C11021 VPWR _489_/a_226_47# 0.12fF
C11022 VPWR _607_/a_78_199# 0.77fF
C11023 _378_/a_558_47# _324_/a_558_47# 0.01fF
C11024 _366_/a_76_199# _366_/a_489_413# 0.12fF
C11025 _328_/A _367_/C 0.23fF
C11026 _378_/A _519_/C 0.10fF
C11027 _418_/B _447_/B 0.02fF
C11028 _371_/B _398_/X 0.11fF
C11029 _596_/a_489_413# VPWR 0.39fF
C11030 _327_/a_78_199# _631_/A 0.19fF
C11031 _375_/X _417_/A 2.88fF
C11032 _410_/B _411_/A 0.05fF
C11033 _461_/a_292_297# _424_/X 0.08fF
C11034 _426_/A _398_/a_489_413# 0.11fF
C11035 _461_/a_78_199# _423_/X 0.15fF
C11036 _390_/B _475_/A 1.02fF
C11037 _330_/A _351_/a_27_53# 0.06fF
C11038 _487_/X _433_/Y 0.05fF
C11039 _614_/a_226_47# M[1] 0.00fF
C11040 _455_/X _356_/a_78_199# 0.17fF
C11041 input10/a_27_47# _397_/a_76_199# 0.01fF
C11042 _530_/a_226_47# _531_/A 0.01fF
C11043 _396_/a_250_297# _392_/A 0.36fF
C11044 _534_/a_209_297# _515_/Y 0.11fF
C11045 VPWR _547_/a_222_93# 0.07fF
C11046 _340_/A _346_/A 0.30fF
C11047 _608_/X _442_/D 0.34fF
C11048 _506_/A _478_/a_27_47# 0.01fF
C11049 _485_/A _410_/C 0.30fF
C11050 _575_/a_215_47# _540_/X 0.03fF
C11051 _575_/a_78_199# _546_/X 0.01fF
C11052 VPWR _591_/A 4.36fF
C11053 _324_/a_62_47# _367_/C 0.45fF
C11054 _393_/A _419_/X 0.03fF
C11055 _510_/X _471_/A 0.01fF
C11056 _597_/a_215_47# _575_/X 0.10fF
C11057 _606_/Y _607_/a_78_199# 0.13fF
C11058 _612_/Y _610_/A 1.28fF
C11059 _623_/X _627_/D 1.54fF
C11060 VPWR _397_/X 1.51fF
C11061 _625_/Y _621_/X 0.26fF
C11062 _627_/C _442_/D 0.03fF
C11063 _454_/X _503_/A 0.07fF
C11064 B[7] _590_/A 0.86fF
C11065 input5/a_381_47# _478_/A 0.69fF
C11066 _519_/X _542_/A 0.17fF
C11067 _380_/A _486_/A 0.19fF
C11068 _433_/Y _438_/X 0.29fF
C11069 _359_/X _359_/B 0.66fF
C11070 _487_/X _540_/X 0.59fF
C11071 _445_/A _631_/A 0.15fF
C11072 VPWR _624_/a_206_369# 0.07fF
C11073 _420_/X _395_/X 0.03fF
C11074 _631_/B _366_/a_489_413# 0.09fF
C11075 _577_/a_489_413# VPWR 0.39fF
C11076 _390_/D _380_/A 0.53fF
C11077 _435_/a_27_47# _570_/B 0.53fF
C11078 _559_/X _616_/A 0.13fF
C11079 _469_/X _472_/B 0.84fF
C11080 A[6] _486_/B 0.28fF
C11081 _389_/a_27_47# _442_/A 0.07fF
C11082 _331_/a_27_47# VPWR 0.58fF
C11083 _404_/a_558_47# _404_/a_841_47# 0.07fF
C11084 _625_/a_27_47# _625_/a_277_47# 0.19fF
C11085 _631_/A _350_/B 0.20fF
C11086 VPWR _518_/X 0.97fF
C11087 _586_/a_76_199# _612_/A 0.24fF
C11088 _567_/Y _530_/X 0.52fF
C11089 _494_/a_226_47# _493_/X 0.57fF
C11090 _623_/a_76_199# M[6] 0.07fF
C11091 _626_/Y _598_/A 0.15fF
C11092 _417_/D _547_/X 0.03fF
C11093 _563_/A _442_/B 0.10fF
C11094 _350_/X _398_/a_76_199# 0.10fF
C11095 _366_/a_226_47# _337_/X 0.57fF
C11096 _471_/A _475_/A 0.07fF
C11097 B[0] _530_/X 0.05fF
C11098 _433_/Y _570_/A 0.15fF
C11099 _516_/a_27_47# _515_/A 0.02fF
C11100 _462_/X _462_/a_76_199# 0.22fF
C11101 _625_/Y _623_/a_226_47# 0.00fF
C11102 _623_/X _623_/a_489_413# 0.01fF
C11103 output25/a_27_47# _442_/B 0.02fF
C11104 _618_/A _625_/a_27_297# 0.19fF
C11105 _356_/a_78_199# _452_/A 0.42fF
C11106 _347_/A _547_/X 0.03fF
C11107 _613_/X M[1] 0.35fF
C11108 _544_/A _486_/X 0.86fF
C11109 _396_/X _392_/A 0.17fF
C11110 _529_/Y _531_/A 0.41fF
C11111 _426_/a_68_297# _426_/A 0.30fF
C11112 _410_/B _334_/a_109_47# 0.02fF
C11113 _456_/a_489_413# _454_/X 0.16fF
C11114 _615_/a_78_199# _573_/A 0.03fF
C11115 _583_/X _582_/Y 0.01fF
C11116 _630_/a_76_199# _629_/X 0.27fF
C11117 _406_/A _631_/Y 0.03fF
C11118 _544_/A _513_/A 0.48fF
C11119 _437_/a_448_47# _437_/X 0.01fF
C11120 _616_/Y _618_/A 1.15fF
C11121 _616_/A _616_/B 1.13fF
C11122 _551_/X _559_/X 0.00fF
C11123 _474_/A _510_/a_68_297# 0.01fF
C11124 _439_/X _468_/X 0.06fF
C11125 _487_/X _378_/A 0.37fF
C11126 _568_/a_227_47# _587_/A 0.04fF
C11127 _418_/a_68_297# _418_/a_150_297# 0.02fF
C11128 _424_/a_76_199# _424_/X 0.22fF
C11129 _540_/X _570_/A 0.04fF
C11130 _487_/X _537_/a_539_297# 0.02fF
C11131 _362_/a_76_199# _351_/X 0.41fF
C11132 _360_/X _436_/A 0.11fF
C11133 _633_/Y _385_/a_558_47# 0.08fF
C11134 _568_/a_539_297# VPWR 0.02fF
C11135 _544_/A _454_/X 0.03fF
C11136 _351_/a_219_297# _351_/X 0.19fF
C11137 _516_/A _381_/B 0.57fF
C11138 _381_/B _539_/A 0.03fF
C11139 _568_/a_77_199# _570_/B 0.19fF
C11140 _417_/D _488_/a_76_199# 0.11fF
C11141 _408_/B _631_/B 0.38fF
C11142 _381_/C _378_/A 0.03fF
C11143 _536_/a_109_297# _547_/X 0.02fF
C11144 _412_/X _458_/a_215_47# 0.12fF
C11145 _396_/a_250_297# _392_/Y 0.03fF
C11146 _396_/a_93_21# _330_/A 0.39fF
C11147 _583_/a_76_199# _581_/B 0.02fF
C11148 _587_/A _510_/A 0.99fF
C11149 _567_/B _493_/a_215_47# 0.16fF
C11150 _520_/X VPWR 8.70fF
C11151 _620_/a_76_199# _618_/A 0.13fF
C11152 _583_/X _613_/X 0.25fF
C11153 _542_/a_109_47# _542_/B 0.01fF
C11154 _542_/C _442_/a_27_47# 0.16fF
C11155 _542_/a_27_47# _542_/C 0.17fF
C11156 _590_/A VPWR 3.82fF
C11157 _437_/a_79_199# VPWR 0.65fF
C11158 _420_/a_448_47# VPWR 0.08fF
C11159 _622_/a_29_53# _622_/a_111_297# 0.01fF
C11160 _351_/X _374_/a_78_199# 0.33fF
C11161 _455_/X _390_/D 0.03fF
C11162 B[2] _577_/a_76_199# 0.18fF
C11163 _469_/A _584_/A 0.22fF
C11164 _611_/a_27_297# _591_/Y 0.24fF
C11165 _397_/X _399_/a_215_47# 0.10fF
C11166 _390_/B _390_/a_197_47# 0.03fF
C11167 _587_/A _485_/D 0.03fF
C11168 _417_/A _337_/B 0.30fF
C11169 VPWR _522_/a_489_413# 0.39fF
C11170 _594_/a_109_297# _593_/Y 0.17fF
C11171 _418_/B _418_/X 0.35fF
C11172 _492_/a_489_413# VPWR 0.39fF
C11173 _630_/a_76_199# _432_/B 0.46fF
C11174 _613_/a_77_199# _586_/a_505_21# 0.00fF
C11175 _533_/X _549_/X 0.56fF
C11176 _563_/A _563_/D 0.34fF
C11177 _608_/a_78_199# _608_/a_292_297# 0.03fF
C11178 _551_/X _550_/X 0.32fF
C11179 _609_/a_209_297# _627_/B 0.01fF
C11180 _506_/Y _511_/a_250_297# 0.00fF
C11181 input5/a_841_47# VPWR 0.31fF
C11182 _375_/X _631_/B 0.03fF
C11183 _473_/a_227_297# _472_/Y 0.03fF
C11184 _523_/a_76_199# _523_/a_489_413# 0.12fF
C11185 _473_/a_77_199# _471_/A 0.17fF
C11186 _473_/a_323_297# _471_/Y 0.01fF
C11187 _318_/a_27_47# VPWR 0.80fF
C11188 _611_/X _627_/C 0.11fF
C11189 VPWR _384_/a_489_413# 0.39fF
C11190 _587_/A _483_/X 0.94fF
C11191 _471_/A _390_/B 1.38fF
C11192 _620_/a_226_47# _620_/a_489_413# 0.02fF
C11193 _620_/a_76_199# _620_/a_226_297# 0.01fF
C11194 _570_/B _588_/A 0.20fF
C11195 _620_/X _606_/A 0.01fF
C11196 _631_/Y _442_/A 0.81fF
C11197 _604_/X _602_/Y 0.29fF
C11198 _532_/a_206_369# _527_/Y 0.15fF
C11199 _532_/a_76_199# _527_/A 0.20fF
X_432_ _432_/A _432_/X _432_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_26_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_501_ _531_/A _501_/Y VGND VPWR _531_/C _531_/A _531_/C VPWR VGND sky130_fd_sc_hd__a2bb2oi_1
X_363_ _363_/A _430_/A _363_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_13_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_13_100 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_346_ VPWR VGND _347_/A _346_/A VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_10_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_415_ VGND VPWR _561_/A _448_/A VPWR VGND sky130_fd_sc_hd__buf_1
X_329_ VGND VPWR VGND VPWR _314_/X _314_/X _328_/X _329_/X _328_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_13 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_9_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_18_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_594_ _573_/A _593_/Y _594_/X _593_/A _573_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__a22o_1
XFILLER_13_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput31 _501_/Y M[8] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_16_120 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput20 _607_/X M[12] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_577_ VGND VPWR VGND VPWR _559_/X _559_/X _576_/X _580_/A _576_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_123 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XTAP_112 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_431_ VGND VPWR VGND VPWR _428_/X _428_/X _430_/X _431_/X _430_/X sky130_fd_sc_hd__a2bb2o_1
X_362_ VGND VPWR VGND VPWR _351_/X _351_/X _361_/X _363_/B _361_/X sky130_fd_sc_hd__a2bb2o_1
X_500_ _464_/A _531_/C _465_/X _427_/A _466_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_3_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_629_ _629_/A _629_/X _629_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_10_148 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_345_ _442_/B _346_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_414_ _542_/A _448_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_328_ _328_/A _328_/X _328_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_9_34 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_593_ _593_/A _593_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_6_13 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_68 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_25_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_15_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_15_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
Xoutput21 _620_/X M[13] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_576_ VGND VPWR VGND VPWR _574_/X _574_/X _575_/X _576_/X _575_/X sky130_fd_sc_hd__a2bb2o_1
Xoutput32 _530_/X M[9] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XTAP_124 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_361_ VGND VPWR VGND VPWR _352_/X _352_/X _360_/X _361_/X _360_/X sky130_fd_sc_hd__a2bb2o_1
X_430_ _430_/A _430_/X _432_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_13_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_9_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_628_ _623_/X _625_/Y _628_/Y _622_/X _621_/X _627_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o221ai_2
XFILLER_3_36 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_559_ _559_/X _535_/Y _570_/A _503_/A _538_/Y _539_/X VPWR VGND VPWR VGND sky130_fd_sc_hd__o32a_1
XFILLER_12_12 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_344_ _338_/X _363_/A _342_/X _329_/X _343_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_413_ _447_/B _413_/X _516_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_23_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_23_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_0_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_3_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_327_ _481_/A _328_/B _367_/C _631_/A _445_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_1_91 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
X_592_ _590_/A _591_/Y _593_/A _590_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__a21oi_1
XFILLER_19_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
Xoutput22 _626_/Y M[14] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_575_ _547_/X _575_/X _540_/X _546_/X _548_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XTAP_125 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ VGND VPWR VGND VPWR _353_/X _353_/X _359_/X _360_/X _359_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_558_ _558_/X _556_/Y _557_/A _557_/B _556_/A _557_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__o32a_1
X_489_ VGND VPWR VGND VPWR _483_/X _483_/X _488_/X _489_/X _488_/X sky130_fd_sc_hd__a2bb2o_1
X_627_ _627_/C _627_/A _627_/X _627_/B _627_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__or4_1
XFILLER_10_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_10_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_7 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_343_ VGND VPWR VGND VPWR _329_/X _329_/X _338_/X _343_/X _338_/X sky130_fd_sc_hd__a2bb2o_1
X_412_ VGND VPWR VGND VPWR _408_/X _408_/X _411_/X _412_/X _411_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_2_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_326_ VGND VPWR _445_/A _326_/A VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_20_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_591_ _591_/A _591_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_15_68 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_15_13 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput23 _628_/Y M[15] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XTAP_126 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_11_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_574_ _572_/B _572_/A _573_/Y _574_/X VPWR VGND VPWR VGND sky130_fd_sc_hd__a21o_1
XFILLER_13_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_557_ _557_/B _557_/Y _557_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
X_626_ _623_/X _626_/Y VGND VPWR _625_/Y _623_/X _625_/Y VPWR VGND sky130_fd_sc_hd__a2bb2oi_1
X_488_ VGND VPWR VGND VPWR _486_/X _486_/X _487_/X _488_/X _487_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_8_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_342_ _350_/C _342_/X _631_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_411_ _411_/A _411_/X _411_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_12_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
X_609_ _469_/X _608_/X _542_/D _622_/C _610_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_23_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_325_ _390_/D _326_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_18_13 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_71 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_590_ _590_/A _591_/A _590_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_19_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_13_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_10_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput24 _633_/Y M[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XTAP_127 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_573_ _573_/A _573_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_22_138 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_7_92 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_26_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_625_ _606_/A _624_/X _625_/Y _601_/A _618_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__a31oi_2
X_556_ _556_/A _556_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_12_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_487_ _452_/X _487_/X _447_/X _449_/A _453_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_341_ VGND VPWR _631_/B _436_/A VPWR VGND sky130_fd_sc_hd__buf_1
X_410_ _411_/B _410_/C _542_/B _410_/B _542_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_10_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_539_ _539_/A _539_/X _587_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_608_ _627_/B _608_/X _627_/C _627_/A _627_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_23_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_324_ VPWR VGND VPWR VGND _448_/B _367_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_20_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_15_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput25 _634_/Y M[2] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_572_ _572_/A _573_/A _572_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XTAP_128 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_60 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_26_47 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_26_36 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_26_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_3_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_3_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_555_ _556_/A _554_/A _554_/X _554_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21bo_1
X_624_ _616_/A _624_/X _616_/B _616_/Y _599_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__o2bb2a_1
X_486_ _486_/A _486_/X _486_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_8_110 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_12_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_340_ _340_/A _350_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_607_ _606_/Y _607_/X _601_/A _601_/Y _606_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_5_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_5_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_146 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_538_ _538_/A _538_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_23_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_469_ VPWR VGND VPWR VGND _469_/A _469_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_105 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_116 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_323_ _417_/A _448_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_1_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_25_159 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_25_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_25_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_15_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xoutput26 _635_/Y M[3] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_16_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_571_ _572_/B _569_/A _570_/X _569_/Y _381_/B _469_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__a32o_1
XTAP_129 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_118 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_21_70 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XTAP_107 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_554_ _554_/A _554_/X _554_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_623_ VGND VPWR VGND VPWR _621_/X _621_/X _622_/X _623_/X _622_/X sky130_fd_sc_hd__a2bb2o_1
X_485_ _486_/B _542_/A _485_/A _542_/D _485_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_399_ _397_/X _426_/A _350_/X _374_/X _398_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_27_91 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_468_ _438_/X _468_/X _436_/X _437_/X _439_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_4_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_606_ _606_/A _606_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_537_ _538_/A _535_/Y _570_/A _472_/B _535_/A _536_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__o32a_1
XFILLER_23_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_322_ _322_/A _481_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_2_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_13_82 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_70 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_20_17 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_72 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
Xoutput27 _373_/Y M[4] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_25_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_127 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_28 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
X_570_ _570_/A _570_/X _570_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XTAP_119 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_13_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_71 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_553_ _524_/X _554_/B _504_/X _523_/X _525_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_12_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_622_ _627_/B _622_/X _627_/D _622_/C VPWR VGND VPWR VGND sky130_fd_sc_hd__or3_1
X_484_ _563_/B _486_/A _561_/A _367_/C _519_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_12_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_398_ VGND VPWR VGND VPWR _374_/X _374_/X _397_/X _398_/X _397_/X sky130_fd_sc_hd__a2bb2o_1
X_467_ _465_/X _467_/Y VGND VPWR _466_/X _465_/X _466_/X VPWR VGND sky130_fd_sc_hd__a2bb2oi_1
X_605_ _602_/Y _604_/X _556_/Y _557_/A _606_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a31o_1
X_536_ _585_/B _536_/Y _570_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
X_321_ _442_/A _322_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_9_19 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_519_ _519_/A _519_/X _563_/B _519_/C VPWR VGND VPWR VGND sky130_fd_sc_hd__or3_1
XFILLER_24_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_24_82 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_10_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xoutput28 _630_/X M[5] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xoutput17 _631_/Y M[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XTAP_109 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_21_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_16_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_552_ VGND VPWR VGND VPWR _533_/X _533_/X _551_/X _554_/A _551_/X sky130_fd_sc_hd__a2bb2o_1
X_483_ _483_/X _480_/Y _480_/A _482_/X _410_/C _386_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__a32o_1
X_621_ _610_/A _621_/X _611_/X _591_/A _613_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_8_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_466_ _430_/X _466_/X _431_/X _428_/X _432_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_397_ VGND VPWR VGND VPWR _384_/X _384_/X _396_/X _397_/X _396_/X sky130_fd_sc_hd__a2bb2o_1
X_604_ _602_/Y _603_/Y _556_/Y _557_/B _604_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a31o_1
X_535_ _535_/A _535_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_23_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_64 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
X_320_ VPWR VGND _631_/A _452_/A VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_13_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_1_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_449_ _449_/A _519_/C VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_518_ _518_/X _515_/Y _515_/A _517_/X _381_/B _386_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__a32o_1
XFILLER_1_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_19_159 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_63 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput18 _558_/X M[10] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_25_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput29 _433_/Y M[6] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_24_162 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_15_140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_21_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_620_ VGND VPWR VGND VPWR _618_/Y _618_/Y _619_/Y _620_/X _619_/Y sky130_fd_sc_hd__a2bb2o_1
X_551_ VGND VPWR VGND VPWR _549_/X _549_/X _550_/X _551_/X _550_/X sky130_fd_sc_hd__a2bb2o_1
X_482_ _539_/A _482_/X _563_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_8_147 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_465_ _427_/A _464_/A _465_/X _464_/Y _427_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__a22o_1
X_396_ _396_/X _392_/Y _392_/A _395_/X _386_/X _330_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__a32o_1
X_603_ VGND VPWR _579_/X _554_/X _581_/B _603_/Y VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_5_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_534_ _386_/A _514_/B _381_/B _515_/Y _535_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_13_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_448_ _448_/A _449_/A _448_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_517_ _570_/A _517_/X _584_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_379_ _516_/A _382_/A _452_/A _448_/B _544_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_1_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_24_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput19 _583_/X M[11] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_15_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XPHY_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_21 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_16_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_8_159 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_481_ VGND VPWR _539_/A _481_/A VPWR VGND sky130_fd_sc_hd__buf_1
X_550_ _521_/X _550_/X _511_/X _520_/X _522_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_27_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_464_ _464_/A _464_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_602_ _602_/A _602_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_533_ _533_/X _506_/Y _539_/A _503_/A _509_/Y _510_/X VPWR VGND VPWR VGND sky130_fd_sc_hd__o32a_1
X_395_ _584_/A _395_/X _436_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_378_ VPWR VGND VPWR VGND _378_/A _544_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_447_ _544_/A _447_/X _447_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_516_ VGND VPWR _570_/A _516_/A VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_24_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_19_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_10_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_21_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_21_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_21_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_16_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_480_ _480_/A _480_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_27_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_601_ _601_/A _601_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_27_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_463_ VGND VPWR VGND VPWR _406_/Y _406_/Y _462_/X _464_/A _462_/X sky130_fd_sc_hd__a2bb2o_1
X_532_ _527_/A _557_/B _527_/B _527_/Y _498_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__o2bb2a_1
X_394_ VPWR VGND VPWR VGND _563_/D _584_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_4_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_446_ _446_/X _444_/Y _444_/A _445_/X _410_/B _386_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__a32o_1
XFILLER_13_21 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_1_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_377_ _380_/A _378_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_515_ _515_/A _515_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_429_ VGND VPWR VGND VPWR _350_/X _350_/X _398_/X _432_/B _398_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xinput1 VGND VPWR _330_/A A[0] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_19_118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XTAP_90 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_86 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_24_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_24_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_21_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XPHY_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_23_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_78 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_531_ _531_/C _557_/A _531_/A _531_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__nor3_1
X_462_ VGND VPWR VGND VPWR _460_/X _460_/X _461_/X _462_/X _461_/X sky130_fd_sc_hd__a2bb2o_1
X_393_ _393_/A _563_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_4_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_4_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_600_ _599_/Y _598_/B _598_/A _601_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_13_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_514_ _514_/A _515_/A _514_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_445_ _445_/A _445_/X _563_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_376_ _447_/B _376_/X _481_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_24_98 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_428_ _426_/B _426_/A _427_/Y _428_/X VPWR VGND VPWR VGND sky130_fd_sc_hd__a21o_1
X_359_ _359_/A _359_/X _359_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
Xinput2 A[1] _390_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XTAP_91 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_56 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XTAP_80 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_152 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_98 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_24_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_24_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_21_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_16_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_15_133 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_21_136 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_12_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_530_ VGND VPWR VGND VPWR _531_/B _531_/B _529_/Y _530_/X _529_/Y sky130_fd_sc_hd__a2bb2o_1
X_461_ _423_/X _461_/X _407_/Y _422_/X _424_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_392_ _392_/A _392_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_4_36 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_47 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_13_89 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_444_ _444_/A _444_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_375_ _359_/B _353_/X _375_/X _359_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ba_1
X_513_ _514_/B _542_/A _513_/A _542_/B _542_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_427_ _427_/A _427_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_358_ _359_/B _381_/C _485_/A _442_/A _381_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_1_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_1_26 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XTAP_92 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 VPWR VGND VPWR VGND A[2] _390_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_81 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_120 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_19_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_24_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_2_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_89 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_8_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_27_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_391_ _391_/A _392_/A _391_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_460_ VGND VPWR VGND VPWR _440_/X _440_/X _459_/X _460_/X _459_/X sky130_fd_sc_hd__a2bb2o_1
X_589_ VGND VPWR VGND VPWR _612_/A _612_/A _588_/Y _590_/B _588_/Y sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_13_13 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_374_ _360_/X _374_/X _351_/X _352_/X _361_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_443_ _443_/A _444_/A _443_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_512_ _347_/A _514_/A _561_/A _378_/A _340_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_24_34 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_426_ _426_/A _427_/A _426_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XTAP_93 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_357_ _478_/A _381_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xinput4 VGND VPWR _442_/A A[3] VPWR VGND sky130_fd_sc_hd__buf_1
XTAP_60 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_67 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_409_ _326_/A _411_/A _481_/A _563_/A _350_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_21_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_2_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_13 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_116 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_105 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_27_45 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_390_ _391_/B _542_/C _542_/B _390_/B _390_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_8_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_588_ _627_/D _588_/Y _588_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
X_373_ _371_/A _629_/B _373_/Y _371_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__a21oi_1
X_442_ _443_/B _478_/A _442_/A _442_/B _442_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_511_ _511_/X _509_/A _510_/X _509_/Y _410_/B _469_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__a32o_1
XFILLER_5_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xinput5 VPWR VGND VPWR VGND A[4] _478_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_425_ VGND VPWR VGND VPWR _407_/Y _407_/Y _424_/X _426_/B _424_/X sky130_fd_sc_hd__a2bb2o_1
X_356_ _481_/A _359_/A _452_/A _448_/B _516_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_27_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_19_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XTAP_94 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ _563_/D _408_/X _408_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_339_ _442_/D _340_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_7_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_14_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_8_92 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_587_ VGND VPWR _627_/D _587_/A VPWR VGND sky130_fd_sc_hd__buf_1
X_372_ _432_/A _629_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_510_ _510_/A _510_/X _587_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_441_ _346_/A _443_/A _355_/A _322_/A _340_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_1_116 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_24_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_424_ VGND VPWR VGND VPWR _422_/X _422_/X _423_/X _424_/X _423_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_355_ VPWR VGND _516_/A _355_/A VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_1_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xinput6 VGND VPWR _380_/A A[5] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_27_101 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XTAP_95 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_49 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XTAP_62 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_24_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_407_ VGND VPWR _406_/B _406_/A _406_/Y _407_/Y VPWR VGND sky130_fd_sc_hd__o21ai_1
X_338_ _337_/A _332_/X _338_/X _337_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ba_1
XFILLER_21_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_15_148 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_11_92 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_16_59 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_7_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_586_ VGND VPWR _586_/S _622_/C _503_/A _612_/A VPWR VGND sky130_fd_sc_hd__mux2_1
X_371_ _371_/A _432_/A _371_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_440_ VGND VPWR VGND VPWR _436_/X _436_/X _439_/X _440_/X _439_/X sky130_fd_sc_hd__a2bb2o_1
X_569_ _569_/A _569_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_24_26 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
X_423_ _383_/X _423_/X _384_/X _375_/X _396_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_354_ _478_/A _355_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_6_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XTAP_96 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 VGND VPWR _542_/A A[6] VPWR VGND sky130_fd_sc_hd__buf_1
XTAP_63 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_406_ _406_/Y _406_/B _406_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nand2_1
X_337_ _337_/A _337_/X _337_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_23_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_21_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xinput10 VGND VPWR _417_/A B[1] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_16_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_14_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_7_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_21_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_4_159 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_585_ _585_/B _622_/C _627_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_1_129 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_370_ _370_/A _371_/B _370_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_499_ _497_/B _497_/A _498_/Y _531_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__a21o_1
X_568_ _569_/A _566_/Y _544_/A _567_/B _566_/A _567_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__o32a_1
X_422_ VGND VPWR VGND VPWR _412_/X _412_/X _421_/X _422_/X _421_/X sky130_fd_sc_hd__a2bb2o_1
X_353_ _519_/A _353_/X _445_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XTAP_97 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 A[7] _542_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XTAP_86 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_405_ _503_/A _406_/B _631_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
X_336_ _510_/A _337_/B _367_/C _631_/A _408_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_18_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_21_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_2_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_11_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_11_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_14_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_319_ _417_/D _452_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
Xinput11 VGND VPWR _485_/D B[2] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_22_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_7_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_17_71 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_584_ _584_/A _590_/A _627_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_12_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_152 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_498_ _498_/A _498_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_567_ _567_/B _567_/Y _588_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
X_421_ VGND VPWR VGND VPWR _419_/X _419_/X _420_/X _421_/X _420_/X sky130_fd_sc_hd__a2bb2o_1
X_352_ _328_/A _314_/X _352_/X _328_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ba_1
XTAP_98 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_619_ VGND VPWR _606_/Y _601_/Y _599_/A _619_/Y VPWR VGND sky130_fd_sc_hd__o21ai_1
XTAP_76 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 VGND VPWR _417_/D B[0] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_27_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_25_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_148 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_335_ VPWR VGND VPWR VGND _445_/A _510_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_404_ VPWR VGND VPWR VGND _585_/B _503_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_21_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_15_118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_11_40 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_318_ _328_/A _485_/A _381_/C _410_/C _390_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
Xinput12 VPWR VGND VPWR VGND B[3] _442_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_22_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_22_72 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_7_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_94 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_583_ VGND VPWR VGND VPWR _602_/A _602_/A _582_/Y _583_/X _582_/Y sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_635_ _635_/Y _370_/A _371_/B _370_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__a21boi_1
X_497_ _497_/A _498_/A _497_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_5_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_566_ _566_/A _566_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_24_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_351_ _351_/A _350_/X _351_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__or2b_1
X_420_ _382_/B _376_/X _420_/X _382_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ba_1
XFILLER_14_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_19_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XTAP_99 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_618_ _618_/A _618_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XTAP_77 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_549_ VGND VPWR VGND VPWR _540_/X _540_/X _548_/X _549_/X _548_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_18_127 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_334_ _337_/A _485_/A _381_/C _410_/B _390_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_403_ VGND VPWR _585_/B _472_/B VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_2_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_98 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_23_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_15_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xinput13 VGND VPWR _442_/B B[4] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_11_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_11_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_317_ VGND VPWR _485_/A _417_/A VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_20_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_11_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_27_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_582_ VGND VPWR _557_/Y _556_/A _554_/X _582_/Y VPWR VGND sky130_fd_sc_hd__o21ai_1
X_496_ _461_/X _497_/B _406_/Y _460_/X _462_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_634_ _634_/Y _368_/A _370_/A _368_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__a21boi_1
XFILLER_0_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
X_565_ _386_/A _543_/B _513_/A _543_/Y _566_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_5_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_98 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_350_ _350_/C _563_/A _350_/X _350_/B _408_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__or4_1
XTAP_89 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_617_ _616_/A _616_/Y _618_/A _616_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__a21oi_1
XTAP_67 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_548_ VGND VPWR VGND VPWR _546_/X _546_/X _547_/X _548_/X _547_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_78 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_479_ _479_/A _480_/A _479_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_27_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_27_128 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_402_ VGND VPWR _472_/B _567_/B VPWR VGND sky130_fd_sc_hd__buf_1
X_333_ VGND VPWR _410_/B _390_/D VPWR VGND sky130_fd_sc_hd__buf_1
Xinput14 VGND VPWR _393_/A B[5] VPWR VGND sky130_fd_sc_hd__buf_1
X_316_ VPWR VGND VPWR VGND _442_/A _410_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_20_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_22_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_27_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_17_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_581_ _602_/A _579_/X _581_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_3_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_495_ VGND VPWR VGND VPWR _468_/X _468_/X _494_/X _497_/A _494_/X sky130_fd_sc_hd__a2bb2o_1
X_633_ _368_/B _633_/Y _633_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2b_1
X_564_ _564_/A _586_/S _572_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_5_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_478_ _479_/B _513_/A _478_/A _542_/B _542_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XTAP_57 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_616_ _616_/B _616_/Y _616_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
X_547_ _486_/B _518_/X _547_/X _519_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ba_1
XTAP_79 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_401_ _401_/A _567_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XPHY_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_332_ _519_/A _332_/X _436_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XPHY_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_2_56 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_45 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_23_143 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_23_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xinput15 VGND VPWR _401_/A B[6] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_20_146 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_315_ VPWR VGND _381_/C _417_/D VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_22_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_11_146 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_135 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_11_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_8_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_580_ _580_/A _581_/B _580_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_632_ _475_/A _633_/A _367_/C _631_/A _631_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_0_145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_563_ _627_/C _563_/A _586_/S _563_/B _563_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__or4_1
X_494_ VGND VPWR VGND VPWR _492_/X _492_/X _493_/X _494_/X _493_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XTAP_58 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_615_ _593_/Y _616_/B _594_/X _573_/A _595_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XTAP_69 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_546_ VGND VPWR VGND VPWR _543_/Y _543_/Y _545_/Y _546_/X _545_/Y sky130_fd_sc_hd__a2bb2o_1
X_477_ _347_/A _479_/A _544_/A _516_/A _340_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_27_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_26_152 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_25_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_331_ VGND VPWR _436_/A _350_/B VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_400_ _330_/A _391_/B _386_/X _392_/Y _406_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a31o_1
XPHY_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_529_ VGND VPWR _531_/C _531_/A _498_/A _529_/Y VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_17_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_17_152 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_23_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_23_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_11_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_11_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_314_ _519_/A _314_/X _408_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_14_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xinput16 VGND VPWR _469_/A B[7] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_20_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_114 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_103 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_22_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_11_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_8_56 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_0_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_90 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_631_ _631_/B _631_/Y _631_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
X_493_ _458_/X _493_/X _440_/X _457_/X _459_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_562_ _627_/B _564_/A _627_/C _563_/A _584_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_5_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_476_ _476_/X _474_/A _475_/X _474_/Y _390_/B _469_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__a32o_1
XFILLER_14_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XTAP_59 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_614_ VGND VPWR VGND VPWR _611_/X _611_/X _613_/X _616_/A _613_/X sky130_fd_sc_hd__a2bb2o_1
X_545_ _584_/A _545_/Y _588_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
XPHY_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_25_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_25_43 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_330_ _330_/A _350_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XPHY_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_459_ VGND VPWR VGND VPWR _457_/X _457_/X _458_/X _459_/X _458_/X sky130_fd_sc_hd__a2bb2o_1
X_528_ _527_/B _527_/A _527_/Y _531_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__a21o_1
XFILLER_11_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_313_ VGND VPWR _408_/B _313_/A VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_14_101 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_26_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_8_68 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_0_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_630_ VGND VPWR VGND VPWR _432_/B _432_/B _629_/X _630_/X _629_/X sky130_fd_sc_hd__a2bb2o_1
X_492_ VGND VPWR VGND VPWR _476_/X _476_/X _491_/X _492_/X _491_/X sky130_fd_sc_hd__a2bb2o_1
X_561_ VGND VPWR _627_/C _561_/A VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_5_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_34 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_14_12 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_613_ _613_/X _612_/Y _588_/A _627_/D _627_/A _586_/S VPWR VGND VPWR VGND sky130_fd_sc_hd__o32a_1
X_475_ _475_/A _475_/X _587_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_544_ VPWR VGND VPWR VGND _544_/A _588_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_26_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_25_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_25_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_458_ _420_/X _458_/X _412_/X _419_/X _421_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_527_ _527_/B _527_/Y _527_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_17_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_389_ VGND VPWR _542_/C _442_/D VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_2_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_312_ _390_/B _313_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_14_146 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_91 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_101 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_3_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_491_ VGND VPWR VGND VPWR _489_/X _489_/X _490_/X _491_/X _490_/X sky130_fd_sc_hd__a2bb2o_1
X_560_ VGND VPWR _627_/B _563_/B VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_5_26 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_68 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_14_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_474_ _474_/A _474_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_612_ _612_/A _612_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_543_ _543_/B _543_/Y _543_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_26_111 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XPHY_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_6_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_25_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_526_ VGND VPWR VGND VPWR _504_/X _504_/X _525_/X _527_/B _525_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_457_ VGND VPWR VGND VPWR _446_/X _446_/X _456_/X _457_/X _456_/X sky130_fd_sc_hd__a2bb2o_1
X_388_ VGND VPWR _542_/B _442_/B VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_14_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_311_ VGND VPWR _519_/A _447_/B VPWR VGND sky130_fd_sc_hd__buf_1
X_509_ _509_/A _509_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_22_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_17_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_490_ _455_/X _490_/X _446_/X _454_/X _456_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_9_91 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_473_ _474_/A _471_/Y _510_/A _472_/B _471_/A _472_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__o32a_1
X_611_ _591_/A _610_/A _611_/X _610_/Y _591_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__a22o_1
X_542_ _543_/B _542_/C _542_/A _542_/B _542_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_25_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_25_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XPHY_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_9_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_387_ _313_/A _391_/A _350_/C _347_/A _445_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_525_ VGND VPWR VGND VPWR _523_/X _523_/X _524_/X _525_/X _524_/X sky130_fd_sc_hd__a2bb2o_1
X_456_ VGND VPWR VGND VPWR _454_/X _454_/X _455_/X _456_/X _455_/X sky130_fd_sc_hd__a2bb2o_1
X_310_ _485_/D _447_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_439_ VGND VPWR VGND VPWR _437_/X _437_/X _438_/X _439_/X _438_/X sky130_fd_sc_hd__a2bb2o_1
X_508_ _509_/A _506_/Y _539_/A _585_/B _506_/A _507_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__o32a_1
XFILLER_8_49 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_147 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_24_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_0_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_0_128 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_472_ _472_/B _472_/Y _510_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
X_610_ _610_/A _610_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_541_ _347_/A _543_/A _340_/A _561_/A _451_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_6_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_524_ _490_/X _524_/X _476_/X _489_/X _491_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_455_ _418_/B _413_/X _455_/X _418_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ba_1
X_386_ VPWR VGND VPWR VGND _386_/A _386_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_369_ VGND VPWR VGND VPWR _342_/X _342_/X _343_/X _370_/B _343_/X sky130_fd_sc_hd__a2bb2o_1
X_438_ _475_/A _438_/X _472_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_507_ _585_/B _507_/Y _539_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_9_120 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_6_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_126 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_471_ _471_/A _471_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
X_540_ _540_/X _538_/A _539_/X _538_/Y _410_/C _469_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__a32o_1
XFILLER_20_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_26_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_26_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_26_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_25_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_136 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_385_ VPWR VGND VPWR VGND _393_/A _386_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_523_ VGND VPWR VGND VPWR _511_/X _511_/X _522_/X _523_/X _522_/X sky130_fd_sc_hd__a2bb2o_1
X_454_ VGND VPWR VGND VPWR _447_/X _447_/X _453_/X _454_/X _453_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_22_150 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_26_91 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_26_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_368_ _368_/A _370_/A _368_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_437_ _411_/B _408_/X _437_/X _411_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ba_1
X_506_ _506_/A _506_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_3_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_146 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_23_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_82 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
X_470_ _386_/A _443_/B _410_/B _444_/Y _471_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a31o_1
X_599_ _599_/A _599_/Y VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_26_148 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_384_ VGND VPWR VGND VPWR _375_/X _375_/X _383_/X _384_/X _383_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_159 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_522_ VGND VPWR VGND VPWR _520_/X _520_/X _521_/X _522_/X _521_/X sky130_fd_sc_hd__a2bb2o_1
X_453_ _453_/X _519_/C _452_/X _449_/A _381_/C _542_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__a32o_1
X_436_ _436_/A _436_/X _587_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_367_ _367_/C _631_/A _368_/B _475_/A _631_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__or4_1
X_505_ _386_/A _479_/B _410_/C _480_/Y _506_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_9_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_26_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_12_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_12_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_6_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__fill_2
XFILLER_17_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_419_ VGND VPWR VGND VPWR _413_/X _413_/X _418_/X _419_/X _418_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_64 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_84 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_50 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_26_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XPHY_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_598_ _598_/A _599_/A _598_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_6_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_25_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XPHY_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_383_ VGND VPWR VGND VPWR _376_/X _376_/X _382_/X _383_/X _382_/X sky130_fd_sc_hd__a2bb2o_1
X_452_ _452_/A _452_/X _563_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_521_ _487_/X _521_/X _483_/X _486_/X _488_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_16_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_61 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XTAP_130 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_22_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_26_71 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_366_ VGND VPWR VGND VPWR _332_/X _332_/X _337_/X _368_/A _337_/X sky130_fd_sc_hd__a2bb2o_1
X_504_ _504_/X _471_/Y _510_/A _627_/A _474_/Y _475_/X VPWR VGND VPWR VGND sky130_fd_sc_hd__o32a_1
XFILLER_13_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_435_ VGND VPWR _587_/A _570_/B VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_9_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_22_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_349_ _436_/A _351_/A _350_/C _563_/A _475_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_418_ _418_/A _418_/X _418_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_23_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_0_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_597_ _575_/X _598_/B _559_/X _574_/X _576_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_6_42 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_520_ VGND VPWR VGND VPWR _518_/X _518_/X _519_/X _520_/X _519_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_382_ _382_/A _382_/X _382_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_1
X_451_ VGND VPWR _563_/B _451_/A VPWR VGND sky130_fd_sc_hd__buf_1
XTAP_120 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_365_ _363_/B _363_/A _629_/A _371_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__a21o_1
X_503_ VPWR VGND VPWR VGND _503_/A _627_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_434_ _469_/A _570_/B VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_9_135 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_3_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_3_43 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_63 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_348_ VGND VPWR _475_/A _408_/B VPWR VGND sky130_fd_sc_hd__buf_1
X_417_ _418_/B _542_/A _417_/A _513_/A _417_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_5_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_119 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_24_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_0_44 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_73 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_20_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_596_ VGND VPWR VGND VPWR _594_/X _594_/X _595_/X _598_/A _595_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_381_ _382_/B _381_/C _485_/A _381_/B _513_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_450_ _542_/D _451_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XTAP_121 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_151 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_579_ VPWR VGND _579_/X _580_/B _580_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_433_ _431_/X _433_/Y VGND VPWR _432_/X _431_/X _432_/X VPWR VGND sky130_fd_sc_hd__a2bb2oi_1
XFILLER_22_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_502_ _493_/X _527_/A _468_/X _492_/X _494_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
X_364_ _430_/A _629_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_13_143 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_22 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_3_66 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_10_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_10_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_12_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_347_ _347_/A _563_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_5_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X_416_ _378_/A _418_/A _561_/A _448_/B _452_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_2_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
XFILLER_9_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_98 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_18_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_18_96 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_595_ _595_/X _566_/Y _588_/A _627_/A _569_/Y _570_/X VPWR VGND VPWR VGND sky130_fd_sc_hd__o32a_1
XFILLER_20_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_25_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
Xoutput30 _467_/Y M[7] VGND VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_17_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_380_ VGND VPWR _513_/A _380_/A VPWR VGND sky130_fd_sc_hd__buf_1
XTAP_122 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X_578_ _550_/X _580_/B _533_/X _549_/X _551_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o22a_1
C11200 _580_/B VGND 1.82fF
C11201 _549_/X VGND 1.70fF
C11202 _578_/a_215_47# VGND 0.68fF **FLOATING
C11203 _578_/a_493_297# VGND 0.00fF **FLOATING
C11204 _578_/a_292_297# VGND 0.00fF **FLOATING
C11205 _578_/a_78_199# VGND 0.52fF **FLOATING
C11206 _380_/a_27_47# VGND 0.69fF **FLOATING
C11207 M[7] VGND 1.29fF
C11208 _467_/Y VGND 0.93fF
C11209 output30/a_27_47# VGND 0.95fF **FLOATING
C11210 _570_/X VGND 1.33fF
C11211 _566_/Y VGND 1.69fF
C11212 _595_/a_227_47# VGND 0.78fF **FLOATING
C11213 _595_/a_77_199# VGND 0.41fF **FLOATING
C11214 _416_/a_215_47# VGND 0.67fF **FLOATING
C11215 _416_/a_78_199# VGND 0.47fF **FLOATING
C11216 _347_/A VGND 4.69fF
C11217 _347_/a_27_47# VGND 0.92fF **FLOATING
C11218 _430_/A VGND 0.75fF
C11219 _502_/a_215_47# VGND 0.67fF **FLOATING
C11220 _502_/a_78_199# VGND 0.45fF **FLOATING
C11221 _433_/a_481_47# VGND 0.01fF **FLOATING
C11222 _433_/a_397_297# VGND 0.06fF **FLOATING
C11223 _433_/a_109_47# VGND 0.85fF **FLOATING
C11224 _579_/X VGND 0.03fF
C11225 _579_/a_59_75# VGND 0.68fF **FLOATING
C11226 _382_/B VGND 3.15fF
C11227 _381_/a_303_47# VGND 0.01fF **FLOATING
C11228 _381_/a_197_47# VGND 0.02fF **FLOATING
C11229 _381_/a_109_47# VGND 0.01fF **FLOATING
C11230 _381_/a_27_47# VGND 0.70fF **FLOATING
C11231 _596_/a_556_47# VGND 0.01fF **FLOATING
C11232 _596_/a_489_413# VGND 0.11fF **FLOATING
C11233 _596_/a_226_47# VGND 0.78fF **FLOATING
C11234 _596_/a_76_199# VGND 0.69fF **FLOATING
C11235 _417_/a_303_47# VGND 0.01fF **FLOATING
C11236 _417_/a_197_47# VGND 0.02fF **FLOATING
C11237 _417_/a_109_47# VGND 0.01fF **FLOATING
C11238 _417_/a_27_47# VGND 0.77fF **FLOATING
C11239 _348_/a_27_47# VGND 0.68fF **FLOATING
C11240 _570_/B VGND 0.60fF
C11241 _469_/A VGND 2.89fF
C11242 _503_/a_841_47# VGND 0.50fF **FLOATING
C11243 _503_/a_664_47# VGND 0.68fF **FLOATING
C11244 _503_/a_558_47# VGND 0.69fF **FLOATING
C11245 _503_/a_381_47# VGND 0.35fF **FLOATING
C11246 _503_/a_62_47# VGND 0.79fF **FLOATING
C11247 _365_/a_384_47# VGND 0.01fF **FLOATING
C11248 _365_/a_299_297# VGND 0.09fF **FLOATING
C11249 _365_/a_81_21# VGND 0.70fF **FLOATING
C11250 _563_/B VGND 4.60fF
C11251 _451_/A VGND 0.77fF
C11252 _451_/a_27_47# VGND 0.69fF **FLOATING
C11253 _382_/a_68_297# VGND 0.53fF **FLOATING
C11254 _520_/a_556_47# VGND 0.01fF **FLOATING
C11255 _520_/a_489_413# VGND 0.10fF **FLOATING
C11256 _520_/a_226_47# VGND 0.81fF **FLOATING
C11257 _520_/a_76_199# VGND 0.70fF **FLOATING
C11258 _598_/B VGND 0.18fF
C11259 _574_/X VGND 2.13fF
C11260 _575_/X VGND 0.14fF
C11261 _576_/X VGND 0.26fF
C11262 _597_/a_215_47# VGND 0.67fF **FLOATING
C11263 _597_/a_78_199# VGND 0.47fF **FLOATING
C11264 _418_/X VGND 1.11fF
C11265 _418_/B VGND 1.05fF
C11266 _418_/a_68_297# VGND 0.55fF **FLOATING
C11267 _351_/A VGND 0.65fF
C11268 _349_/a_215_47# VGND 0.58fF **FLOATING
C11269 _349_/a_78_199# VGND 0.47fF **FLOATING
C11270 _435_/a_27_47# VGND 0.69fF **FLOATING
C11271 _504_/a_227_47# VGND 0.80fF **FLOATING
C11272 _504_/a_77_199# VGND 0.39fF **FLOATING
C11273 _337_/X VGND 2.34fF
C11274 _366_/a_556_47# VGND 0.01fF **FLOATING
C11275 _366_/a_226_297# VGND 0.00fF **FLOATING
C11276 _366_/a_489_413# VGND 0.17fF **FLOATING
C11277 _366_/a_226_47# VGND 0.63fF **FLOATING
C11278 _366_/a_76_199# VGND 0.24fF **FLOATING
C11279 _521_/a_215_47# VGND 0.67fF **FLOATING
C11280 _521_/a_493_297# VGND 0.00fF **FLOATING
C11281 _521_/a_292_297# VGND 0.00fF **FLOATING
C11282 _452_/X VGND 2.09fF
C11283 _452_/a_68_297# VGND 0.55fF **FLOATING
C11284 _383_/X VGND 4.32fF
C11285 _383_/a_556_47# VGND 0.01fF **FLOATING
C11286 _383_/a_489_413# VGND 0.11fF **FLOATING
C11287 _383_/a_226_47# VGND 0.77fF **FLOATING
C11288 _383_/a_76_199# VGND 0.71fF **FLOATING
C11289 _598_/a_68_297# VGND 0.53fF **FLOATING
C11290 _419_/a_556_47# VGND 0.01fF **FLOATING
C11291 _419_/a_489_413# VGND 0.10fF **FLOATING
C11292 _419_/a_226_47# VGND 0.81fF **FLOATING
C11293 _419_/a_76_199# VGND 0.70fF **FLOATING
C11294 _505_/a_303_47# VGND 0.01fF **FLOATING
C11295 _505_/a_209_47# VGND 0.01fF **FLOATING
C11296 _505_/a_209_297# VGND 0.03fF **FLOATING
C11297 _505_/a_80_21# VGND 0.74fF **FLOATING
C11298 _367_/a_27_297# VGND 0.94fF **FLOATING
C11299 _436_/a_68_297# VGND 0.54fF **FLOATING
C11300 _453_/a_584_47# VGND 0.01fF **FLOATING
C11301 _453_/a_346_47# VGND 0.02fF **FLOATING
C11302 _453_/a_256_47# VGND 0.01fF **FLOATING
C11303 _453_/a_250_297# VGND 0.05fF **FLOATING
C11304 _453_/a_93_21# VGND 0.77fF **FLOATING
C11305 _521_/X VGND 0.38fF
C11306 _522_/a_556_47# VGND 0.01fF **FLOATING
C11307 _522_/a_489_413# VGND 0.10fF **FLOATING
C11308 _522_/a_226_47# VGND 0.77fF **FLOATING
C11309 _522_/a_76_199# VGND 0.67fF **FLOATING
C11310 _384_/a_556_47# VGND 0.01fF **FLOATING
C11311 _384_/a_489_413# VGND 0.11fF **FLOATING
C11312 _384_/a_226_47# VGND 0.75fF **FLOATING
C11313 _384_/a_76_199# VGND 0.70fF **FLOATING
C11314 _470_/a_303_47# VGND 0.01fF **FLOATING
C11315 _470_/a_209_47# VGND 0.01fF **FLOATING
C11316 _470_/a_209_297# VGND 0.03fF **FLOATING
C11317 _470_/a_80_21# VGND 0.72fF **FLOATING
C11318 _506_/Y VGND 0.07fF
C11319 _506_/A VGND 0.43fF
C11320 _408_/X VGND 0.22fF
C11321 _437_/a_448_47# VGND 0.42fF **FLOATING
C11322 _437_/a_544_297# VGND 0.01fF **FLOATING
C11323 _437_/a_222_93# VGND 0.55fF **FLOATING
C11324 _437_/a_79_199# VGND 0.69fF **FLOATING
C11325 _368_/a_68_297# VGND 0.55fF **FLOATING
C11326 _453_/X VGND 3.22fF
C11327 _447_/X VGND 4.38fF
C11328 _454_/a_556_47# VGND 0.01fF **FLOATING
C11329 _454_/a_489_413# VGND 0.10fF **FLOATING
C11330 _454_/a_226_47# VGND 0.79fF **FLOATING
C11331 _454_/a_76_199# VGND 0.70fF **FLOATING
C11332 _523_/X VGND 1.43fF
C11333 _523_/a_556_47# VGND 0.01fF **FLOATING
C11334 _523_/a_489_413# VGND 0.11fF **FLOATING
C11335 _523_/a_226_47# VGND 0.79fF **FLOATING
C11336 _523_/a_76_199# VGND 0.70fF **FLOATING
C11337 _393_/A VGND 4.62fF
C11338 _385_/a_841_47# VGND 0.42fF **FLOATING
C11339 _385_/a_664_47# VGND 0.66fF **FLOATING
C11340 _385_/a_558_47# VGND 0.68fF **FLOATING
C11341 _385_/a_381_47# VGND 0.35fF **FLOATING
C11342 _385_/a_62_47# VGND 0.85fF **FLOATING
C11343 _410_/C VGND 7.37fF
C11344 _540_/a_584_47# VGND 0.01fF **FLOATING
C11345 _540_/a_346_47# VGND 0.02fF **FLOATING
C11346 _540_/a_256_47# VGND 0.01fF **FLOATING
C11347 _540_/a_250_297# VGND 0.10fF **FLOATING
C11348 _540_/a_93_21# VGND 0.88fF **FLOATING
C11349 _438_/X VGND 1.72fF
C11350 _438_/a_68_297# VGND 0.55fF **FLOATING
C11351 _370_/B VGND 0.51fF
C11352 _369_/a_556_47# VGND 0.01fF **FLOATING
C11353 _369_/a_489_413# VGND 0.10fF **FLOATING
C11354 _369_/a_226_47# VGND 0.76fF **FLOATING
C11355 _369_/a_76_199# VGND 0.71fF **FLOATING
C11356 _386_/X VGND 0.62fF
C11357 _386_/a_841_47# VGND 0.50fF **FLOATING
C11358 _386_/a_664_47# VGND 0.68fF **FLOATING
C11359 _386_/a_558_47# VGND 0.70fF **FLOATING
C11360 _386_/a_381_47# VGND 0.36fF **FLOATING
C11361 _386_/a_62_47# VGND 0.81fF **FLOATING
C11362 _413_/X VGND 2.44fF
C11363 _455_/a_448_47# VGND 0.53fF **FLOATING
C11364 _455_/a_222_93# VGND 0.46fF **FLOATING
C11365 _455_/a_79_199# VGND 0.55fF **FLOATING
C11366 _490_/X VGND 1.35fF
C11367 _491_/X VGND 1.46fF
C11368 _476_/X VGND 3.24fF
C11369 _524_/a_215_47# VGND 0.66fF **FLOATING
C11370 _524_/a_78_199# VGND 0.41fF **FLOATING
C11371 _340_/A VGND 3.26fF
C11372 _541_/a_215_47# VGND 0.58fF **FLOATING
C11373 _541_/a_78_199# VGND 0.38fF **FLOATING
C11374 _610_/Y VGND 0.51fF
C11375 _472_/a_109_297# VGND 0.04fF **FLOATING
C11376 _509_/A VGND 1.80fF
C11377 _508_/a_227_47# VGND 0.80fF **FLOATING
C11378 _508_/a_77_199# VGND 0.39fF **FLOATING
C11379 _439_/a_556_47# VGND 0.01fF **FLOATING
C11380 _439_/a_489_413# VGND 0.10fF **FLOATING
C11381 _439_/a_226_47# VGND 0.81fF **FLOATING
C11382 _439_/a_76_199# VGND 0.71fF **FLOATING
C11383 _447_/B VGND 3.29fF
C11384 _456_/X VGND 3.58fF
C11385 _456_/a_556_47# VGND 0.01fF **FLOATING
C11386 _456_/a_489_413# VGND 0.11fF **FLOATING
C11387 _456_/a_226_47# VGND 0.70fF **FLOATING
C11388 _456_/a_76_199# VGND 0.71fF **FLOATING
C11389 _525_/a_556_47# VGND 0.01fF **FLOATING
C11390 _525_/a_489_413# VGND 0.10fF **FLOATING
C11391 _525_/a_226_47# VGND 0.77fF **FLOATING
C11392 _525_/a_76_199# VGND 0.67fF **FLOATING
C11393 _391_/A VGND 1.52fF
C11394 _313_/A VGND 1.87fF
C11395 _387_/a_215_47# VGND 0.60fF **FLOATING
C11396 _387_/a_78_199# VGND 0.47fF **FLOATING
C11397 _542_/C VGND 7.16fF
C11398 _542_/a_303_47# VGND 0.01fF **FLOATING
C11399 _542_/a_197_47# VGND 0.02fF **FLOATING
C11400 _542_/a_109_47# VGND 0.01fF **FLOATING
C11401 _542_/a_27_47# VGND 0.69fF **FLOATING
C11402 _611_/a_373_47# VGND 0.01fF **FLOATING
C11403 _611_/a_109_47# VGND 0.04fF **FLOATING
C11404 _611_/a_109_297# VGND 0.07fF **FLOATING
C11405 _611_/a_27_297# VGND 1.09fF **FLOATING
C11406 _471_/A VGND 2.14fF
C11407 _472_/Y VGND 0.54fF
C11408 _473_/a_227_47# VGND 0.81fF **FLOATING
C11409 _473_/a_77_199# VGND 0.39fF **FLOATING
C11410 _446_/X VGND 0.54fF
C11411 _490_/a_215_47# VGND 0.67fF **FLOATING
C11412 _490_/a_78_199# VGND 0.43fF **FLOATING
C11413 _509_/Y VGND 0.84fF
C11414 _519_/A VGND 7.06fF
C11415 _311_/a_27_47# VGND 0.66fF **FLOATING
C11416 _388_/a_27_47# VGND 0.66fF **FLOATING
C11417 _457_/X VGND 3.42fF
C11418 _457_/a_556_47# VGND 0.01fF **FLOATING
C11419 _457_/a_489_413# VGND 0.11fF **FLOATING
C11420 _457_/a_226_47# VGND 0.70fF **FLOATING
C11421 _457_/a_76_199# VGND 0.71fF **FLOATING
C11422 _527_/B VGND 1.55fF
C11423 _526_/a_556_47# VGND 0.01fF **FLOATING
C11424 _526_/a_489_413# VGND 0.11fF **FLOATING
C11425 _526_/a_226_47# VGND 0.79fF **FLOATING
C11426 _526_/a_76_199# VGND 0.68fF **FLOATING
C11427 _543_/Y VGND 1.18fF
C11428 _474_/Y VGND 2.61fF
C11429 _474_/A VGND 0.75fF
C11430 _560_/a_27_47# VGND 0.66fF **FLOATING
C11431 _491_/a_556_47# VGND 0.01fF **FLOATING
C11432 _491_/a_489_413# VGND 0.10fF **FLOATING
C11433 _491_/a_226_47# VGND 0.78fF **FLOATING
C11434 _491_/a_76_199# VGND 0.70fF **FLOATING
C11435 _389_/a_27_47# VGND 0.67fF **FLOATING
C11436 _421_/X VGND 1.44fF
C11437 _458_/a_215_47# VGND 0.67fF **FLOATING
C11438 _458_/a_78_199# VGND 0.44fF **FLOATING
C11439 _544_/a_841_47# VGND 0.50fF **FLOATING
C11440 _544_/a_664_47# VGND 0.67fF **FLOATING
C11441 _544_/a_558_47# VGND 0.68fF **FLOATING
C11442 _544_/a_381_47# VGND 0.35fF **FLOATING
C11443 _544_/a_62_47# VGND 0.79fF **FLOATING
C11444 _475_/A VGND 0.81fF
C11445 _475_/a_68_297# VGND 0.56fF **FLOATING
C11446 _627_/A VGND 1.06fF
C11447 _586_/S VGND 1.51fF
C11448 _612_/Y VGND 5.62fF
C11449 _613_/a_227_47# VGND 0.80fF **FLOATING
C11450 _613_/a_77_199# VGND 0.40fF **FLOATING
C11451 _627_/C VGND 7.20fF
C11452 _561_/A VGND 0.92fF
C11453 _561_/a_27_47# VGND 0.66fF **FLOATING
C11454 _492_/a_556_47# VGND 0.01fF **FLOATING
C11455 _492_/a_489_413# VGND 0.11fF **FLOATING
C11456 _492_/a_226_47# VGND 0.75fF **FLOATING
C11457 _492_/a_76_199# VGND 0.69fF **FLOATING
C11458 _630_/X VGND 2.00fF
C11459 _629_/X VGND 0.06fF
C11460 _630_/a_556_47# VGND 0.01fF **FLOATING
C11461 _630_/a_489_413# VGND 0.10fF **FLOATING
C11462 _630_/a_226_47# VGND 0.77fF **FLOATING
C11463 _630_/a_76_199# VGND 0.71fF **FLOATING
C11464 _313_/a_27_47# VGND 0.77fF **FLOATING
C11465 _527_/A VGND 1.28fF
C11466 _527_/Y VGND 1.51fF
C11467 _528_/a_384_47# VGND 0.01fF **FLOATING
C11468 _528_/a_299_297# VGND 0.09fF **FLOATING
C11469 _528_/a_81_21# VGND 0.70fF **FLOATING
C11470 _458_/X VGND 0.46fF
C11471 _459_/X VGND 1.73fF
C11472 _459_/a_556_47# VGND 0.01fF **FLOATING
C11473 _459_/a_489_413# VGND 0.10fF **FLOATING
C11474 _459_/a_226_47# VGND 0.71fF **FLOATING
C11475 _459_/a_76_199# VGND 0.72fF **FLOATING
C11476 _611_/X VGND 0.87fF
C11477 _614_/a_556_47# VGND 0.01fF **FLOATING
C11478 _614_/a_489_413# VGND 0.10fF **FLOATING
C11479 _614_/a_226_47# VGND 0.68fF **FLOATING
C11480 _614_/a_76_199# VGND 0.69fF **FLOATING
C11481 _475_/X VGND 0.65fF
C11482 _476_/a_584_47# VGND 0.01fF **FLOATING
C11483 _476_/a_346_47# VGND 0.02fF **FLOATING
C11484 _476_/a_256_47# VGND 0.01fF **FLOATING
C11485 _476_/a_250_297# VGND 0.03fF **FLOATING
C11486 _476_/a_93_21# VGND 0.64fF **FLOATING
C11487 _563_/A VGND 6.70fF
C11488 _562_/a_215_47# VGND 0.58fF **FLOATING
C11489 _562_/a_292_297# VGND 0.00fF **FLOATING
C11490 _493_/a_215_47# VGND 0.68fF **FLOATING
C11491 _493_/a_78_199# VGND 0.42fF **FLOATING
C11492 B[7] VGND 9.88fF
C11493 input16/a_27_47# VGND 0.72fF **FLOATING
C11494 _314_/X VGND 0.74fF
C11495 _314_/a_68_297# VGND 0.54fF **FLOATING
C11496 _529_/a_27_47# VGND 0.47fF **FLOATING
C11497 _330_/A VGND 1.99fF
C11498 _400_/a_303_47# VGND 0.03fF **FLOATING
C11499 _400_/a_209_47# VGND 0.01fF **FLOATING
C11500 _400_/a_209_297# VGND 0.10fF **FLOATING
C11501 _400_/a_80_21# VGND 0.32fF **FLOATING
C11502 _331_/a_27_47# VGND 0.67fF **FLOATING
C11503 _477_/a_215_47# VGND 0.67fF **FLOATING
C11504 _477_/a_493_297# VGND 0.00fF **FLOATING
C11505 _477_/a_292_297# VGND 0.00fF **FLOATING
C11506 _477_/a_78_199# VGND 0.51fF **FLOATING
C11507 _546_/a_556_47# VGND 0.01fF **FLOATING
C11508 _546_/a_489_413# VGND 0.11fF **FLOATING
C11509 _546_/a_226_47# VGND 0.78fF **FLOATING
C11510 _546_/a_76_199# VGND 0.70fF **FLOATING
C11511 _595_/X VGND 0.96fF
C11512 _594_/X VGND 1.08fF
C11513 _615_/a_215_47# VGND 0.68fF **FLOATING
C11514 _615_/a_78_199# VGND 0.45fF **FLOATING
C11515 _494_/a_556_47# VGND 0.01fF **FLOATING
C11516 _494_/a_489_413# VGND 0.11fF **FLOATING
C11517 _494_/a_226_47# VGND 0.81fF **FLOATING
C11518 _494_/a_76_199# VGND 0.70fF **FLOATING
C11519 _563_/D VGND 7.03fF
C11520 _563_/a_27_297# VGND 0.93fF **FLOATING
C11521 _633_/A VGND 0.65fF
C11522 _632_/a_215_47# VGND 0.56fF **FLOATING
C11523 _632_/a_78_199# VGND 0.47fF **FLOATING
C11524 _581_/B VGND 0.51fF
C11525 _580_/a_68_297# VGND 0.56fF **FLOATING
C11526 _417_/D VGND 2.63fF
C11527 _315_/a_161_47# VGND 1.10fF **FLOATING
C11528 B[6] VGND 1.24fF
C11529 input15/a_75_212# VGND 0.67fF **FLOATING
C11530 _332_/X VGND 3.88fF
C11531 _332_/a_150_297# VGND 0.00fF **FLOATING
C11532 _332_/a_68_297# VGND 0.66fF **FLOATING
C11533 _401_/A VGND 1.23fF
C11534 _547_/a_448_47# VGND 0.50fF **FLOATING
C11535 _547_/a_222_93# VGND 0.46fF **FLOATING
C11536 _547_/a_79_199# VGND 0.54fF **FLOATING
C11537 _478_/a_303_47# VGND 0.01fF **FLOATING
C11538 _478_/a_197_47# VGND 0.02fF **FLOATING
C11539 _478_/a_109_47# VGND 0.01fF **FLOATING
C11540 _478_/a_27_47# VGND 0.75fF **FLOATING
C11541 _564_/A VGND 1.53fF
C11542 _564_/a_27_53# VGND 0.80fF **FLOATING
C11543 _564_/a_219_297# VGND 0.58fF **FLOATING
C11544 _368_/B VGND 2.20fF
C11545 _633_/a_74_47# VGND 0.56fF **FLOATING
C11546 _494_/X VGND 1.29fF
C11547 _468_/X VGND 1.74fF
C11548 _495_/a_556_47# VGND 0.01fF **FLOATING
C11549 _495_/a_489_413# VGND 0.12fF **FLOATING
C11550 _495_/a_226_47# VGND 0.79fF **FLOATING
C11551 _495_/a_76_199# VGND 0.70fF **FLOATING
C11552 _581_/a_206_47# VGND 0.01fF **FLOATING
C11553 _581_/a_27_93# VGND 0.59fF **FLOATING
C11554 _316_/a_841_47# VGND 0.55fF **FLOATING
C11555 _316_/a_664_47# VGND 0.66fF **FLOATING
C11556 _316_/a_558_47# VGND 0.69fF **FLOATING
C11557 _316_/a_381_47# VGND 0.37fF **FLOATING
C11558 _316_/a_62_47# VGND 0.80fF **FLOATING
C11559 B[5] VGND 2.47fF
C11560 _333_/a_27_47# VGND 0.69fF **FLOATING
C11561 _402_/a_27_47# VGND 0.78fF **FLOATING
C11562 _479_/A VGND 1.20fF
C11563 _479_/B VGND 1.27fF
C11564 _479_/a_68_297# VGND 0.63fF **FLOATING
C11565 _548_/a_556_47# VGND 0.01fF **FLOATING
C11566 _548_/a_489_413# VGND 0.10fF **FLOATING
C11567 _548_/a_226_47# VGND 0.76fF **FLOATING
C11568 _548_/a_76_199# VGND 0.67fF **FLOATING
C11569 _616_/B VGND 2.98fF
C11570 _616_/A VGND 0.80fF
C11571 _616_/Y VGND 1.03fF
C11572 _617_/a_199_47# VGND 0.01fF **FLOATING
C11573 _617_/a_113_297# VGND 0.09fF **FLOATING
C11574 _350_/X VGND 3.11fF
C11575 _350_/B VGND 1.09fF
C11576 _350_/a_277_297# VGND 0.00fF **FLOATING
C11577 _350_/a_205_297# VGND 0.00fF **FLOATING
C11578 _350_/a_109_297# VGND 0.00fF **FLOATING
C11579 _350_/a_27_297# VGND 0.91fF **FLOATING
C11580 _565_/a_303_47# VGND 0.01fF **FLOATING
C11581 _565_/a_80_21# VGND 0.70fF **FLOATING
C11582 _634_/Y VGND 2.13fF
C11583 _634_/a_384_47# VGND 0.01fF **FLOATING
C11584 _634_/a_300_297# VGND 0.03fF **FLOATING
C11585 _634_/a_27_413# VGND 0.70fF **FLOATING
C11586 _461_/X VGND 2.95fF
C11587 _462_/X VGND 0.80fF
C11588 _406_/Y VGND 3.29fF
C11589 _496_/a_215_47# VGND 0.67fF **FLOATING
C11590 _496_/a_78_199# VGND 0.43fF **FLOATING
C11591 _557_/Y VGND 1.59fF
C11592 _582_/a_27_47# VGND 0.46fF **FLOATING
C11593 _317_/a_27_47# VGND 0.73fF **FLOATING
C11594 B[4] VGND 1.37fF
C11595 input13/a_27_47# VGND 0.64fF **FLOATING
C11596 _403_/a_27_47# VGND 0.77fF **FLOATING
C11597 _337_/A VGND 2.85fF
C11598 _390_/B VGND 1.68fF
C11599 _334_/a_303_47# VGND 0.01fF **FLOATING
C11600 _334_/a_197_47# VGND 0.02fF **FLOATING
C11601 _334_/a_109_47# VGND 0.01fF **FLOATING
C11602 _334_/a_27_47# VGND 0.70fF **FLOATING
C11603 _549_/a_556_47# VGND 0.01fF **FLOATING
C11604 _549_/a_489_413# VGND 0.11fF **FLOATING
C11605 _549_/a_226_47# VGND 0.80fF **FLOATING
C11606 _549_/a_76_199# VGND 0.69fF **FLOATING
C11607 _420_/a_448_47# VGND 0.53fF **FLOATING
C11608 _420_/a_222_93# VGND 0.49fF **FLOATING
C11609 _420_/a_79_199# VGND 0.55fF **FLOATING
C11610 _351_/X VGND 1.42fF
C11611 _351_/a_27_53# VGND 0.79fF **FLOATING
C11612 _351_/a_219_297# VGND 0.63fF **FLOATING
C11613 _497_/a_68_297# VGND 0.54fF **FLOATING
C11614 _635_/Y VGND 0.61fF
C11615 _635_/a_384_47# VGND 0.01fF **FLOATING
C11616 _635_/a_300_297# VGND 0.03fF **FLOATING
C11617 _635_/a_27_413# VGND 0.81fF **FLOATING
C11618 _583_/a_556_47# VGND 0.01fF **FLOATING
C11619 _583_/a_489_413# VGND 0.11fF **FLOATING
C11620 _583_/a_226_47# VGND 0.79fF **FLOATING
C11621 _583_/a_76_199# VGND 0.69fF **FLOATING
C11622 _442_/D VGND 8.19fF
C11623 B[3] VGND 1.27fF
C11624 input12/a_841_47# VGND 0.50fF **FLOATING
C11625 input12/a_664_47# VGND 0.68fF **FLOATING
C11626 input12/a_558_47# VGND 0.69fF **FLOATING
C11627 input12/a_381_47# VGND 0.36fF **FLOATING
C11628 input12/a_62_47# VGND 0.85fF **FLOATING
C11629 _328_/A VGND 3.51fF
C11630 _318_/a_303_47# VGND 0.01fF **FLOATING
C11631 _318_/a_197_47# VGND 0.02fF **FLOATING
C11632 _318_/a_109_47# VGND 0.01fF **FLOATING
C11633 _318_/a_27_47# VGND 0.74fF **FLOATING
C11634 _404_/a_841_47# VGND 0.55fF **FLOATING
C11635 _404_/a_664_47# VGND 0.69fF **FLOATING
C11636 _404_/a_558_47# VGND 0.70fF **FLOATING
C11637 _404_/a_381_47# VGND 0.35fF **FLOATING
C11638 _404_/a_62_47# VGND 0.81fF **FLOATING
C11639 _335_/a_841_47# VGND 0.49fF **FLOATING
C11640 _335_/a_664_47# VGND 0.68fF **FLOATING
C11641 _335_/a_558_47# VGND 0.71fF **FLOATING
C11642 _335_/a_381_47# VGND 0.38fF **FLOATING
C11643 _335_/a_62_47# VGND 0.81fF **FLOATING
C11644 B[0] VGND 5.11fF
C11645 input9/a_27_47# VGND 0.76fF **FLOATING
C11646 _599_/A VGND 1.26fF
C11647 _606_/Y VGND 0.50fF
C11648 _619_/a_27_47# VGND 0.46fF **FLOATING
C11649 _352_/X VGND 2.09fF
C11650 _352_/a_448_47# VGND 0.50fF **FLOATING
C11651 _352_/a_222_93# VGND 0.46fF **FLOATING
C11652 _352_/a_79_199# VGND 0.53fF **FLOATING
C11653 _421_/a_556_47# VGND 0.01fF **FLOATING
C11654 _421_/a_489_413# VGND 0.11fF **FLOATING
C11655 _421_/a_226_47# VGND 0.80fF **FLOATING
C11656 _421_/a_76_199# VGND 0.69fF **FLOATING
C11657 _584_/a_68_297# VGND 0.57fF **FLOATING
C11658 input11/a_27_47# VGND 0.70fF **FLOATING
C11659 _337_/B VGND 0.90fF
C11660 _336_/a_215_47# VGND 0.79fF **FLOATING
C11661 _336_/a_493_297# VGND 0.01fF **FLOATING
C11662 _336_/a_292_297# VGND 0.01fF **FLOATING
C11663 _336_/a_78_199# VGND 0.67fF **FLOATING
C11664 input8/a_27_47# VGND 0.95fF **FLOATING
C11665 _445_/A VGND 4.05fF
C11666 _353_/a_68_297# VGND 0.58fF **FLOATING
C11667 _422_/a_556_47# VGND 0.01fF **FLOATING
C11668 _422_/a_489_413# VGND 0.10fF **FLOATING
C11669 _422_/a_226_47# VGND 0.80fF **FLOATING
C11670 _422_/a_76_199# VGND 0.69fF **FLOATING
C11671 _566_/A VGND 4.22fF
C11672 _567_/Y VGND 1.05fF
C11673 _568_/a_227_47# VGND 0.80fF **FLOATING
C11674 _568_/a_77_199# VGND 0.41fF **FLOATING
C11675 _497_/B VGND 0.31fF
C11676 _499_/a_384_47# VGND 0.01fF **FLOATING
C11677 _499_/a_299_297# VGND 0.09fF **FLOATING
C11678 _499_/a_81_21# VGND 0.71fF **FLOATING
C11679 _370_/a_68_297# VGND 0.53fF **FLOATING
C11680 _585_/B VGND 12.08fF
C11681 input10/a_27_47# VGND 0.68fF **FLOATING
C11682 _337_/a_68_297# VGND 0.57fF **FLOATING
C11683 _406_/a_113_47# VGND 0.01fF **FLOATING
C11684 A[6] VGND 3.49fF
C11685 input7/a_27_47# VGND 0.66fF **FLOATING
C11686 _423_/a_215_47# VGND 0.67fF **FLOATING
C11687 _423_/a_78_199# VGND 0.41fF **FLOATING
C11688 _439_/X VGND 0.40fF
C11689 _440_/X VGND 2.35fF
C11690 _440_/a_556_47# VGND 0.01fF **FLOATING
C11691 _440_/a_489_413# VGND 0.10fF **FLOATING
C11692 _440_/a_226_47# VGND 0.79fF **FLOATING
C11693 _440_/a_76_199# VGND 0.69fF **FLOATING
C11694 _432_/A VGND 1.61fF
C11695 _371_/a_68_297# VGND 0.56fF **FLOATING
C11696 _586_/a_439_47# VGND 0.01fF **FLOATING
C11697 _586_/a_218_47# VGND 0.01fF **FLOATING
C11698 _586_/a_505_21# VGND 0.71fF **FLOATING
C11699 _586_/a_76_199# VGND 0.67fF **FLOATING
C11700 _338_/X VGND 1.22fF
C11701 _338_/a_448_47# VGND 0.50fF **FLOATING
C11702 _338_/a_222_93# VGND 0.47fF **FLOATING
C11703 _338_/a_79_199# VGND 0.54fF **FLOATING
C11704 _407_/Y VGND 1.22fF
C11705 _407_/a_27_47# VGND 0.45fF **FLOATING
C11706 A[5] VGND 2.30fF
C11707 input6/a_27_47# VGND 0.66fF **FLOATING
C11708 _355_/a_161_47# VGND 1.11fF **FLOATING
C11709 _424_/a_556_47# VGND 0.01fF **FLOATING
C11710 _424_/a_489_413# VGND 0.11fF **FLOATING
C11711 _424_/a_226_47# VGND 0.77fF **FLOATING
C11712 _424_/a_76_199# VGND 0.69fF **FLOATING
C11713 _441_/a_215_47# VGND 0.58fF **FLOATING
C11714 _441_/a_292_297# VGND 0.00fF **FLOATING
C11715 _510_/A VGND 1.72fF
C11716 _510_/a_68_297# VGND 0.54fF **FLOATING
C11717 _587_/a_27_47# VGND 0.63fF **FLOATING
C11718 _408_/a_68_297# VGND 0.56fF **FLOATING
C11719 _359_/A VGND 1.95fF
C11720 _356_/a_215_47# VGND 0.67fF **FLOATING
C11721 _356_/a_78_199# VGND 0.43fF **FLOATING
C11722 _426_/B VGND 1.11fF
C11723 _425_/a_556_47# VGND 0.01fF **FLOATING
C11724 _425_/a_489_413# VGND 0.10fF **FLOATING
C11725 _425_/a_226_47# VGND 0.80fF **FLOATING
C11726 _425_/a_76_199# VGND 0.69fF **FLOATING
C11727 A[4] VGND 1.84fF
C11728 input5/a_841_47# VGND 0.49fF **FLOATING
C11729 input5/a_664_47# VGND 0.66fF **FLOATING
C11730 input5/a_558_47# VGND 0.69fF **FLOATING
C11731 input5/a_381_47# VGND 0.35fF **FLOATING
C11732 input5/a_62_47# VGND 0.90fF **FLOATING
C11733 _410_/B VGND 6.63fF
C11734 _511_/a_584_47# VGND 0.01fF **FLOATING
C11735 _511_/a_346_47# VGND 0.02fF **FLOATING
C11736 _511_/a_256_47# VGND 0.01fF **FLOATING
C11737 _511_/a_250_297# VGND 0.05fF **FLOATING
C11738 _511_/a_93_21# VGND 0.79fF **FLOATING
C11739 _442_/a_303_47# VGND 0.01fF **FLOATING
C11740 _442_/a_197_47# VGND 0.02fF **FLOATING
C11741 _442_/a_109_47# VGND 0.01fF **FLOATING
C11742 _442_/a_27_47# VGND 0.74fF **FLOATING
C11743 _373_/a_199_47# VGND 0.01fF **FLOATING
C11744 _373_/a_113_297# VGND 0.09fF **FLOATING
C11745 _588_/Y VGND 1.12fF
C11746 _588_/A VGND 6.75fF
C11747 _391_/B VGND 1.49fF
C11748 _390_/a_303_47# VGND 0.01fF **FLOATING
C11749 _390_/a_197_47# VGND 0.02fF **FLOATING
C11750 _390_/a_109_47# VGND 0.01fF **FLOATING
C11751 _390_/a_27_47# VGND 0.75fF **FLOATING
C11752 _326_/A VGND 1.08fF
C11753 _409_/a_215_47# VGND 0.67fF **FLOATING
C11754 _409_/a_78_199# VGND 0.42fF **FLOATING
C11755 _442_/A VGND 5.19fF
C11756 A[3] VGND 3.60fF
C11757 input4/a_27_47# VGND 0.78fF **FLOATING
C11758 _357_/a_27_47# VGND 0.72fF **FLOATING
C11759 _426_/A VGND 3.82fF
C11760 _426_/a_68_297# VGND 0.58fF **FLOATING
C11761 _512_/a_215_47# VGND 0.67fF **FLOATING
C11762 _512_/a_78_199# VGND 0.43fF **FLOATING
C11763 _443_/a_68_297# VGND 0.56fF **FLOATING
C11764 _374_/a_215_47# VGND 0.70fF **FLOATING
C11765 _374_/a_78_199# VGND 0.49fF **FLOATING
C11766 _612_/A VGND 1.61fF
C11767 _589_/a_556_47# VGND 0.01fF **FLOATING
C11768 _589_/a_489_413# VGND 0.10fF **FLOATING
C11769 _589_/a_226_47# VGND 0.78fF **FLOATING
C11770 _589_/a_76_199# VGND 0.55fF **FLOATING
C11771 _460_/X VGND 1.20fF
C11772 _460_/a_556_47# VGND 0.01fF **FLOATING
C11773 _460_/a_489_413# VGND 0.11fF **FLOATING
C11774 _460_/a_226_47# VGND 0.77fF **FLOATING
C11775 _460_/a_76_199# VGND 0.68fF **FLOATING
C11776 _391_/a_68_297# VGND 0.56fF **FLOATING
C11777 _390_/D VGND 5.54fF
C11778 A[2] VGND 1.23fF
C11779 input3/a_841_47# VGND 0.49fF **FLOATING
C11780 input3/a_664_47# VGND 0.66fF **FLOATING
C11781 input3/a_558_47# VGND 0.69fF **FLOATING
C11782 input3/a_381_47# VGND 0.38fF **FLOATING
C11783 input3/a_62_47# VGND 0.85fF **FLOATING
C11784 _359_/B VGND 2.31fF
C11785 _358_/a_303_47# VGND 0.01fF **FLOATING
C11786 _358_/a_197_47# VGND 0.02fF **FLOATING
C11787 _358_/a_109_47# VGND 0.01fF **FLOATING
C11788 _358_/a_27_47# VGND 0.74fF **FLOATING
C11789 _427_/Y VGND 1.19fF
C11790 _513_/A VGND 1.85fF
C11791 _513_/a_303_47# VGND 0.01fF **FLOATING
C11792 _513_/a_197_47# VGND 0.02fF **FLOATING
C11793 _513_/a_109_47# VGND 0.01fF **FLOATING
C11794 _513_/a_27_47# VGND 0.76fF **FLOATING
C11795 _375_/X VGND 3.72fF
C11796 _375_/a_448_47# VGND 0.50fF **FLOATING
C11797 _375_/a_222_93# VGND 0.50fF **FLOATING
C11798 _375_/a_79_199# VGND 0.53fF **FLOATING
C11799 _422_/X VGND 0.90fF
C11800 _423_/X VGND 3.98fF
C11801 _424_/X VGND 1.65fF
C11802 _461_/a_215_47# VGND 0.67fF **FLOATING
C11803 _461_/a_78_199# VGND 0.43fF **FLOATING
C11804 _529_/Y VGND 2.03fF
C11805 _530_/a_556_47# VGND 0.01fF **FLOATING
C11806 _530_/a_489_413# VGND 0.11fF **FLOATING
C11807 _530_/a_226_47# VGND 0.79fF **FLOATING
C11808 _530_/a_76_199# VGND 0.72fF **FLOATING
C11809 A[1] VGND 0.84fF
C11810 input2/a_27_47# VGND 0.89fF **FLOATING
C11811 _359_/X VGND 2.10fF
C11812 _359_/a_68_297# VGND 0.54fF **FLOATING
C11813 _428_/a_384_47# VGND 0.01fF **FLOATING
C11814 _428_/a_299_297# VGND 0.09fF **FLOATING
C11815 _428_/a_81_21# VGND 0.85fF **FLOATING
C11816 _376_/X VGND 1.48fF
C11817 _376_/a_68_297# VGND 0.55fF **FLOATING
C11818 _445_/a_68_297# VGND 0.56fF **FLOATING
C11819 _515_/A VGND 0.46fF
C11820 _514_/B VGND 1.97fF
C11821 _514_/a_68_297# VGND 0.54fF **FLOATING
C11822 _598_/A VGND 0.95fF
C11823 _600_/a_285_47# VGND 0.01fF **FLOATING
C11824 _600_/a_114_47# VGND 0.01fF **FLOATING
C11825 _600_/a_27_297# VGND 0.13fF **FLOATING
C11826 _462_/a_556_47# VGND 0.01fF **FLOATING
C11827 _462_/a_489_413# VGND 0.11fF **FLOATING
C11828 _462_/a_226_47# VGND 0.80fF **FLOATING
C11829 _462_/a_76_199# VGND 0.73fF **FLOATING
C11830 A[0] VGND 1.97fF
C11831 input1/a_27_47# VGND 0.66fF **FLOATING
C11832 _398_/X VGND 2.10fF
C11833 _429_/a_556_47# VGND 0.01fF **FLOATING
C11834 _429_/a_489_413# VGND 0.10fF **FLOATING
C11835 _429_/a_226_47# VGND 0.80fF **FLOATING
C11836 _429_/a_76_199# VGND 0.68fF **FLOATING
C11837 _515_/Y VGND 0.47fF
C11838 _378_/A VGND 6.86fF
C11839 _445_/X VGND 1.03fF
C11840 _446_/a_584_47# VGND 0.01fF **FLOATING
C11841 _446_/a_346_47# VGND 0.02fF **FLOATING
C11842 _446_/a_256_47# VGND 0.01fF **FLOATING
C11843 _446_/a_250_297# VGND 0.03fF **FLOATING
C11844 _446_/a_93_21# VGND 0.77fF **FLOATING
C11845 _394_/a_841_47# VGND 0.48fF **FLOATING
C11846 _394_/a_664_47# VGND 0.77fF **FLOATING
C11847 _394_/a_558_47# VGND 0.78fF **FLOATING
C11848 _394_/a_381_47# VGND 0.47fF **FLOATING
C11849 _394_/a_62_47# VGND 0.47fF **FLOATING
C11850 _532_/a_489_47# VGND 0.52fF **FLOATING
C11851 _532_/a_205_47# VGND 0.01fF **FLOATING
C11852 _532_/a_206_369# VGND 0.60fF **FLOATING
C11853 _532_/a_76_199# VGND 0.48fF **FLOATING
C11854 _463_/a_556_47# VGND 0.01fF **FLOATING
C11855 _463_/a_489_413# VGND 0.10fF **FLOATING
C11856 _463_/a_226_47# VGND 0.78fF **FLOATING
C11857 _463_/a_76_199# VGND 0.70fF **FLOATING
C11858 _480_/Y VGND 0.98fF
C11859 _480_/A VGND 1.89fF
C11860 _516_/a_27_47# VGND 0.68fF **FLOATING
C11861 _447_/a_68_297# VGND 0.55fF **FLOATING
C11862 _378_/a_841_47# VGND 0.49fF **FLOATING
C11863 _378_/a_664_47# VGND 0.67fF **FLOATING
C11864 _378_/a_558_47# VGND 0.70fF **FLOATING
C11865 _378_/a_381_47# VGND 0.35fF **FLOATING
C11866 _378_/a_62_47# VGND 0.70fF **FLOATING
C11867 _395_/X VGND 0.83fF
C11868 _395_/a_68_297# VGND 0.55fF **FLOATING
C11869 _533_/a_227_47# VGND 0.81fF **FLOATING
C11870 _533_/a_77_199# VGND 0.38fF **FLOATING
C11871 _602_/Y VGND 0.91fF
C11872 _464_/Y VGND 2.04fF
C11873 _511_/X VGND 0.45fF
C11874 _550_/a_215_47# VGND 0.67fF **FLOATING
C11875 _550_/a_78_199# VGND 0.44fF **FLOATING
C11876 _539_/A VGND 0.98fF
C11877 _481_/a_27_47# VGND 0.73fF **FLOATING
C11878 M[11] VGND 1.28fF
C11879 output19/a_27_47# VGND 0.95fF **FLOATING
C11880 _382_/A VGND 1.04fF
C11881 _379_/a_215_47# VGND 0.58fF **FLOATING
C11882 _379_/a_493_297# VGND 0.00fF **FLOATING
C11883 _379_/a_292_297# VGND 0.00fF **FLOATING
C11884 _379_/a_78_199# VGND 0.56fF **FLOATING
C11885 _517_/a_150_297# VGND 0.00fF **FLOATING
C11886 _517_/a_68_297# VGND 0.13fF **FLOATING
C11887 _448_/B VGND 1.98fF
C11888 _448_/a_68_297# VGND 0.54fF **FLOATING
C11889 _534_/a_303_47# VGND 0.01fF **FLOATING
C11890 _534_/a_209_47# VGND 0.01fF **FLOATING
C11891 _534_/a_209_297# VGND 0.02fF **FLOATING
C11892 _534_/a_80_21# VGND 0.75fF **FLOATING
C11893 _603_/Y VGND 1.22fF
C11894 _554_/X VGND 4.87fF
C11895 _603_/a_27_47# VGND 0.42fF **FLOATING
C11896 _396_/X VGND 0.27fF
C11897 _396_/a_584_47# VGND 0.01fF **FLOATING
C11898 _396_/a_346_47# VGND 0.02fF **FLOATING
C11899 _396_/a_256_47# VGND 0.01fF **FLOATING
C11900 _396_/a_250_297# VGND 0.03fF **FLOATING
C11901 _396_/a_93_21# VGND 0.78fF **FLOATING
C11902 _465_/a_373_47# VGND 0.01fF **FLOATING
C11903 _465_/a_109_47# VGND 0.04fF **FLOATING
C11904 _465_/a_109_297# VGND 0.07fF **FLOATING
C11905 _465_/a_27_297# VGND 0.98fF **FLOATING
C11906 _482_/a_68_297# VGND 0.56fF **FLOATING
C11907 _551_/a_556_47# VGND 0.01fF **FLOATING
C11908 _551_/a_489_413# VGND 0.10fF **FLOATING
C11909 _551_/a_226_47# VGND 0.78fF **FLOATING
C11910 _551_/a_76_199# VGND 0.67fF **FLOATING
C11911 _620_/X VGND 0.10fF
C11912 _620_/a_556_47# VGND 0.01fF **FLOATING
C11913 _620_/a_489_413# VGND 0.10fF **FLOATING
C11914 _620_/a_226_47# VGND 0.77fF **FLOATING
C11915 _620_/a_76_199# VGND 0.70fF **FLOATING
C11916 M[6] VGND 5.16fF
C11917 _433_/Y VGND 0.95fF
C11918 output29/a_27_47# VGND 0.98fF **FLOATING
C11919 M[10] VGND 3.61fF
C11920 output18/a_27_47# VGND 0.94fF **FLOATING
C11921 _518_/X VGND 1.46fF
C11922 _518_/a_584_47# VGND 0.02fF **FLOATING
C11923 _518_/a_346_47# VGND 0.02fF **FLOATING
C11924 _518_/a_256_47# VGND 0.01fF **FLOATING
C11925 _518_/a_93_21# VGND 0.63fF **FLOATING
C11926 _449_/A VGND 0.93fF
C11927 _320_/a_161_47# VGND 1.10fF **FLOATING
C11928 _557_/B VGND 0.20fF
C11929 _604_/a_303_47# VGND 0.01fF **FLOATING
C11930 _604_/a_209_47# VGND 0.01fF **FLOATING
C11931 _604_/a_209_297# VGND 0.02fF **FLOATING
C11932 _604_/a_80_21# VGND 0.72fF **FLOATING
C11933 _397_/X VGND 0.91fF
C11934 _397_/a_556_47# VGND 0.01fF **FLOATING
C11935 _397_/a_489_413# VGND 0.10fF **FLOATING
C11936 _397_/a_226_47# VGND 0.77fF **FLOATING
C11937 _397_/a_76_199# VGND 0.72fF **FLOATING
C11938 _428_/X VGND 1.37fF
C11939 _430_/X VGND 1.13fF
C11940 _432_/X VGND 1.70fF
C11941 _431_/X VGND 1.64fF
C11942 _466_/a_215_47# VGND 0.66fF **FLOATING
C11943 _466_/a_78_199# VGND 0.45fF **FLOATING
C11944 _621_/X VGND 4.36fF
C11945 _591_/A VGND 1.76fF
C11946 _621_/a_215_47# VGND 0.75fF **FLOATING
C11947 _621_/a_78_199# VGND 0.47fF **FLOATING
C11948 _483_/a_584_47# VGND 0.01fF **FLOATING
C11949 _483_/a_346_47# VGND 0.02fF **FLOATING
C11950 _483_/a_256_47# VGND 0.01fF **FLOATING
C11951 _483_/a_250_297# VGND 0.04fF **FLOATING
C11952 _483_/a_93_21# VGND 0.78fF **FLOATING
C11953 _552_/a_556_47# VGND 0.01fF **FLOATING
C11954 _552_/a_489_413# VGND 0.10fF **FLOATING
C11955 _552_/a_226_47# VGND 0.77fF **FLOATING
C11956 _552_/a_76_199# VGND 0.69fF **FLOATING
C11957 M[0] VGND 1.49fF
C11958 _631_/Y VGND 1.39fF
C11959 output17/a_27_47# VGND 0.94fF **FLOATING
C11960 M[5] VGND 3.09fF
C11961 output28/a_27_47# VGND 0.84fF **FLOATING
C11962 _519_/X VGND 0.79fF
C11963 _519_/a_29_53# VGND 0.95fF **FLOATING
C11964 _322_/A VGND 1.86fF
C11965 _536_/Y VGND 0.79fF
C11966 _604_/X VGND 0.00fF
C11967 _605_/a_303_47# VGND 0.01fF **FLOATING
C11968 _605_/a_209_47# VGND 0.01fF **FLOATING
C11969 _605_/a_209_297# VGND 0.02fF **FLOATING
C11970 _605_/a_80_21# VGND 0.73fF **FLOATING
C11971 _467_/a_481_47# VGND 0.01fF **FLOATING
C11972 _467_/a_397_297# VGND 0.07fF **FLOATING
C11973 _467_/a_109_47# VGND 0.83fF **FLOATING
C11974 _398_/a_556_47# VGND 0.01fF **FLOATING
C11975 _398_/a_489_413# VGND 0.10fF **FLOATING
C11976 _398_/a_226_47# VGND 0.76fF **FLOATING
C11977 _398_/a_76_199# VGND 0.67fF **FLOATING
C11978 _486_/A VGND 0.70fF
C11979 _367_/C VGND 5.36fF
C11980 _484_/a_215_47# VGND 0.67fF **FLOATING
C11981 _484_/a_78_199# VGND 0.44fF **FLOATING
C11982 _627_/B VGND 1.86fF
C11983 _622_/C VGND 2.88fF
C11984 _622_/a_29_53# VGND 0.98fF **FLOATING
C11985 _553_/a_215_47# VGND 0.67fF **FLOATING
C11986 _553_/a_78_199# VGND 0.46fF **FLOATING
C11987 _570_/A VGND 0.04fF
C11988 _570_/a_68_297# VGND 0.55fF **FLOATING
C11989 M[4] VGND 1.39fF
C11990 output27/a_27_47# VGND 1.02fF **FLOATING
C11991 _322_/a_27_47# VGND 0.89fF **FLOATING
C11992 _472_/B VGND 1.85fF
C11993 _537_/a_227_47# VGND 0.81fF **FLOATING
C11994 _537_/a_77_199# VGND 0.41fF **FLOATING
C11995 _437_/X VGND 2.17fF
C11996 _436_/X VGND 2.47fF
C11997 _468_/a_215_47# VGND 0.76fF **FLOATING
C11998 _468_/a_493_297# VGND 0.01fF **FLOATING
C11999 _468_/a_292_297# VGND 0.01fF **FLOATING
C12000 _468_/a_78_199# VGND 0.60fF **FLOATING
C12001 _399_/a_215_47# VGND 0.67fF **FLOATING
C12002 _399_/a_78_199# VGND 0.43fF **FLOATING
C12003 _486_/B VGND 0.72fF
C12004 _485_/a_303_47# VGND 0.01fF **FLOATING
C12005 _485_/a_197_47# VGND 0.02fF **FLOATING
C12006 _485_/a_109_47# VGND 0.01fF **FLOATING
C12007 _485_/a_27_47# VGND 0.72fF **FLOATING
C12008 _623_/a_556_47# VGND 0.01fF **FLOATING
C12009 _623_/a_489_413# VGND 0.10fF **FLOATING
C12010 _623_/a_226_47# VGND 0.77fF **FLOATING
C12011 _623_/a_76_199# VGND 0.68fF **FLOATING
C12012 _554_/a_68_297# VGND 0.56fF **FLOATING
C12013 _571_/a_584_47# VGND 0.01fF **FLOATING
C12014 _571_/a_346_47# VGND 0.01fF **FLOATING
C12015 _571_/a_256_47# VGND 0.01fF **FLOATING
C12016 _571_/a_250_297# VGND 0.03fF **FLOATING
C12017 _571_/a_93_21# VGND 0.78fF **FLOATING
C12018 output26/a_27_47# VGND 0.91fF **FLOATING
C12019 _469_/a_841_47# VGND 0.51fF **FLOATING
C12020 _469_/a_664_47# VGND 0.67fF **FLOATING
C12021 _469_/a_558_47# VGND 0.69fF **FLOATING
C12022 _469_/a_381_47# VGND 0.36fF **FLOATING
C12023 _469_/a_62_47# VGND 0.80fF **FLOATING
C12024 _538_/Y VGND 2.10fF
C12025 _538_/A VGND 1.45fF
C12026 _607_/a_215_47# VGND 0.68fF **FLOATING
C12027 _607_/a_78_199# VGND 0.47fF **FLOATING
C12028 _350_/C VGND 0.37fF
C12029 _340_/a_27_47# VGND 0.80fF **FLOATING
C12030 _486_/a_68_297# VGND 0.58fF **FLOATING
C12031 _624_/a_489_47# VGND 0.49fF **FLOATING
C12032 _624_/a_205_47# VGND 0.01fF **FLOATING
C12033 _624_/a_206_369# VGND 0.59fF **FLOATING
C12034 _624_/a_76_199# VGND 0.48fF **FLOATING
C12035 _556_/A VGND 2.22fF
C12036 _555_/a_382_47# VGND 0.01fF **FLOATING
C12037 _555_/a_298_297# VGND 0.02fF **FLOATING
C12038 _555_/a_215_297# VGND 0.94fF **FLOATING
C12039 _555_/a_27_413# VGND 0.72fF **FLOATING
C12040 VPWR VGND 752.46fF
C12041 _572_/a_150_297# VGND 0.02fF **FLOATING
C12042 _572_/a_68_297# VGND 0.66fF **FLOATING
C12043 output25/a_27_47# VGND 0.85fF **FLOATING
C12044 _324_/a_841_47# VGND 0.50fF **FLOATING
C12045 _324_/a_664_47# VGND 0.67fF **FLOATING
C12046 _324_/a_558_47# VGND 0.69fF **FLOATING
C12047 _324_/a_381_47# VGND 0.36fF **FLOATING
C12048 _324_/a_62_47# VGND 0.79fF **FLOATING
C12049 _608_/X VGND 0.43fF
C12050 _608_/a_215_47# VGND 0.70fF **FLOATING
C12051 _608_/a_78_199# VGND 0.47fF **FLOATING
C12052 _539_/a_68_297# VGND 0.58fF **FLOATING
C12053 _411_/B VGND 2.26fF
C12054 _410_/a_303_47# VGND 0.01fF **FLOATING
C12055 _410_/a_197_47# VGND 0.02fF **FLOATING
C12056 _410_/a_109_47# VGND 0.01fF **FLOATING
C12057 _410_/a_27_47# VGND 0.74fF **FLOATING
C12058 _436_/A VGND 4.78fF
C12059 _341_/a_27_47# VGND 0.68fF **FLOATING
C12060 _487_/a_215_47# VGND 0.67fF **FLOATING
C12061 _487_/a_78_199# VGND 0.46fF **FLOATING
C12062 _624_/X VGND 1.03fF
C12063 _601_/A VGND 1.88fF
C12064 _606_/A VGND 0.70fF
C12065 _625_/a_277_47# VGND 0.35fF **FLOATING
C12066 _625_/a_27_47# VGND 0.28fF **FLOATING
C12067 _625_/a_27_297# VGND 0.08fF **FLOATING
C12068 _573_/Y VGND 0.48fF
C12069 _573_/A VGND 1.91fF
C12070 M[1] VGND 1.37fF
C12071 output24/a_27_47# VGND 0.71fF **FLOATING
C12072 _590_/a_68_297# VGND 0.58fF **FLOATING
C12073 _542_/D VGND 2.23fF
C12074 _609_/a_303_47# VGND 0.01fF **FLOATING
C12075 _609_/a_209_47# VGND 0.01fF **FLOATING
C12076 _609_/a_209_297# VGND 0.02fF **FLOATING
C12077 _609_/a_80_21# VGND 0.73fF **FLOATING
C12078 _411_/X VGND 2.47fF
C12079 _411_/a_68_297# VGND 0.55fF **FLOATING
C12080 _342_/X VGND 3.14fF
C12081 _342_/a_68_297# VGND 0.57fF **FLOATING
C12082 _488_/a_556_47# VGND 0.01fF **FLOATING
C12083 _488_/a_226_297# VGND 0.00fF **FLOATING
C12084 _488_/a_489_413# VGND 0.05fF **FLOATING
C12085 _488_/a_226_47# VGND 0.85fF **FLOATING
C12086 _488_/a_76_199# VGND 0.80fF **FLOATING
C12087 _625_/Y VGND 3.59fF
C12088 _626_/a_481_47# VGND 0.01fF **FLOATING
C12089 _626_/a_397_297# VGND 0.06fF **FLOATING
C12090 _626_/a_109_47# VGND 0.82fF **FLOATING
C12091 _574_/a_384_47# VGND 0.01fF **FLOATING
C12092 _574_/a_299_297# VGND 0.10fF **FLOATING
C12093 _574_/a_81_21# VGND 0.71fF **FLOATING
C12094 output23/a_27_47# VGND 0.89fF **FLOATING
C12095 _591_/Y VGND 0.83fF
C12096 _326_/a_27_47# VGND 0.69fF **FLOATING
C12097 _412_/X VGND 1.86fF
C12098 _412_/a_556_47# VGND 0.01fF **FLOATING
C12099 _412_/a_489_413# VGND 0.11fF **FLOATING
C12100 _412_/a_226_47# VGND 0.78fF **FLOATING
C12101 _412_/a_76_199# VGND 0.68fF **FLOATING
C12102 _343_/a_556_47# VGND 0.01fF **FLOATING
C12103 _343_/a_489_413# VGND 0.10fF **FLOATING
C12104 _343_/a_226_47# VGND 0.77fF **FLOATING
C12105 _343_/a_76_199# VGND 0.72fF **FLOATING
C12106 _627_/a_27_297# VGND 0.95fF **FLOATING
C12107 _489_/X VGND 1.93fF
C12108 _489_/a_556_47# VGND 0.01fF **FLOATING
C12109 _489_/a_489_413# VGND 0.11fF **FLOATING
C12110 _489_/a_226_47# VGND 0.69fF **FLOATING
C12111 _489_/a_76_199# VGND 0.71fF **FLOATING
C12112 _558_/a_227_47# VGND 0.90fF **FLOATING
C12113 _558_/a_539_297# VGND 0.02fF **FLOATING
C12114 _558_/a_323_297# VGND 0.02fF **FLOATING
C12115 _558_/a_227_297# VGND 0.01fF **FLOATING
C12116 _558_/a_77_199# VGND 0.59fF **FLOATING
C12117 _353_/X VGND 1.08fF
C12118 _360_/X VGND 2.32fF
C12119 _360_/a_556_47# VGND 0.01fF **FLOATING
C12120 _360_/a_489_413# VGND 0.10fF **FLOATING
C12121 _360_/a_226_47# VGND 0.78fF **FLOATING
C12122 _360_/a_76_199# VGND 0.70fF **FLOATING
C12123 _546_/X VGND 0.89fF
C12124 _548_/X VGND 0.51fF
C12125 _575_/a_215_47# VGND 0.67fF **FLOATING
C12126 _575_/a_78_199# VGND 0.45fF **FLOATING
C12127 M[14] VGND 1.16fF
C12128 output22/a_27_47# VGND 0.95fF **FLOATING
C12129 _592_/a_199_47# VGND 0.01fF **FLOATING
C12130 _592_/a_113_297# VGND 0.08fF **FLOATING
C12131 _328_/B VGND 1.96fF
C12132 _327_/a_215_47# VGND 0.58fF **FLOATING
C12133 _327_/a_78_199# VGND 0.46fF **FLOATING
C12134 _413_/a_68_297# VGND 0.54fF **FLOATING
C12135 _329_/X VGND 1.82fF
C12136 _343_/X VGND 2.19fF
C12137 _344_/a_215_47# VGND 0.66fF **FLOATING
C12138 _344_/a_78_199# VGND 0.44fF **FLOATING
C12139 _559_/a_227_47# VGND 0.80fF **FLOATING
C12140 _559_/a_77_199# VGND 0.41fF **FLOATING
C12141 _628_/a_300_47# VGND 1.18fF **FLOATING
C12142 _628_/a_28_47# VGND 0.57fF **FLOATING
C12143 _628_/a_734_297# VGND 0.02fF **FLOATING
C12144 _432_/B VGND 2.52fF
C12145 _430_/a_68_297# VGND 0.53fF **FLOATING
C12146 _361_/X VGND 2.89fF
C12147 _361_/a_556_47# VGND 0.01fF **FLOATING
C12148 _361_/a_489_413# VGND 0.11fF **FLOATING
C12149 _361_/a_226_47# VGND 0.77fF **FLOATING
C12150 _361_/a_76_199# VGND 0.69fF **FLOATING
C12151 output32/a_27_47# VGND 0.88fF **FLOATING
C12152 _576_/a_556_47# VGND 0.01fF **FLOATING
C12153 _576_/a_489_413# VGND 0.11fF **FLOATING
C12154 _576_/a_226_47# VGND 0.76fF **FLOATING
C12155 _576_/a_76_199# VGND 0.67fF **FLOATING
C12156 M[13] VGND 1.59fF
C12157 output21/a_27_47# VGND 0.94fF **FLOATING
C12158 _328_/a_68_297# VGND 0.56fF **FLOATING
C12159 _346_/A VGND 0.31fF
C12160 _629_/a_68_297# VGND 0.54fF **FLOATING
C12161 _427_/A VGND 3.23fF
C12162 _465_/X VGND 2.09fF
C12163 _500_/a_215_47# VGND 0.69fF **FLOATING
C12164 _500_/a_78_199# VGND 0.45fF **FLOATING
C12165 _362_/a_556_47# VGND 0.01fF **FLOATING
C12166 _362_/a_489_413# VGND 0.11fF **FLOATING
C12167 _362_/a_226_47# VGND 0.80fF **FLOATING
C12168 _362_/a_76_199# VGND 0.68fF **FLOATING
C12169 _431_/a_556_47# VGND 0.01fF **FLOATING
C12170 _431_/a_489_413# VGND 0.10fF **FLOATING
C12171 _431_/a_226_47# VGND 0.77fF **FLOATING
C12172 _431_/a_76_199# VGND 0.73fF **FLOATING
C12173 _580_/A VGND 2.33fF
C12174 _577_/a_556_47# VGND 0.01fF **FLOATING
C12175 _577_/a_489_413# VGND 0.12fF **FLOATING
C12176 _577_/a_226_47# VGND 0.79fF **FLOATING
C12177 _577_/a_76_199# VGND 0.68fF **FLOATING
C12178 M[12] VGND 1.82fF
C12179 _607_/X VGND 2.43fF
C12180 output20/a_27_47# VGND 0.96fF **FLOATING
C12181 M[8] VGND 3.27fF
C12182 output31/a_27_47# VGND 0.94fF **FLOATING
C12183 _594_/a_373_47# VGND 0.01fF **FLOATING
C12184 _594_/a_109_47# VGND 0.04fF **FLOATING
C12185 _594_/a_109_297# VGND 0.07fF **FLOATING
C12186 _594_/a_27_297# VGND 0.98fF **FLOATING
C12187 _329_/a_556_47# VGND 0.01fF **FLOATING
C12188 _329_/a_489_413# VGND 0.11fF **FLOATING
C12189 _329_/a_226_47# VGND 0.79fF **FLOATING
C12190 _329_/a_76_199# VGND 0.69fF **FLOATING
C12191 _448_/A VGND 0.46fF
C12192 _415_/a_27_47# VGND 0.64fF **FLOATING
C12193 _346_/a_161_47# VGND 1.09fF **FLOATING
C12194 _363_/A VGND 6.08fF
C12195 _363_/B VGND 2.33fF
C12196 _363_/a_68_297# VGND 0.56fF **FLOATING
C12197 _501_/a_481_47# VGND 0.01fF **FLOATING
C12198 _501_/a_397_297# VGND 0.06fF **FLOATING
C12199 _501_/a_109_47# VGND 0.83fF **FLOATING
C12200 _432_/a_68_297# VGND 0.53fF **FLOATING
// .ends

.option scale = 10000u


.tran 1ns 20ns

.control 
run
.endc
.ends

magic
tech sky130A
magscale 1 2
timestamp 1629484537
<< obsli1 >>
rect 1104 2159 16715 17425
<< obsm1 >>
rect 14 1980 17558 17456
<< metal2 >>
rect 18 18928 74 19728
rect 2042 18928 2098 19728
rect 4066 18928 4122 19728
rect 5906 18928 5962 19728
rect 7930 18928 7986 19728
rect 9770 18928 9826 19728
rect 11794 18928 11850 19728
rect 13634 18928 13690 19728
rect 15658 18928 15714 19728
rect 17498 18928 17554 19728
rect 18 0 74 800
rect 1858 0 1914 800
rect 3882 0 3938 800
rect 5722 0 5778 800
rect 7746 0 7802 800
rect 9586 0 9642 800
rect 11610 0 11666 800
rect 13450 0 13506 800
rect 15474 0 15530 800
rect 17498 0 17554 800
<< obsm2 >>
rect 130 18872 1986 18928
rect 2154 18872 4010 18928
rect 4178 18872 5850 18928
rect 6018 18872 7874 18928
rect 8042 18872 9714 18928
rect 9882 18872 11738 18928
rect 11906 18872 13578 18928
rect 13746 18872 15602 18928
rect 15770 18872 17442 18928
rect 20 856 17552 18872
rect 130 734 1802 856
rect 1970 734 3826 856
rect 3994 734 5666 856
rect 5834 734 7690 856
rect 7858 734 9530 856
rect 9698 734 11554 856
rect 11722 734 13394 856
rect 13562 734 15418 856
rect 15586 734 17442 856
<< metal3 >>
rect 0 17144 800 17264
rect 16784 16872 17584 16992
rect 0 14152 800 14272
rect 16784 13880 17584 14000
rect 0 11432 800 11552
rect 16784 11160 17584 11280
rect 0 8440 800 8560
rect 16784 8168 17584 8288
rect 0 5720 800 5840
rect 16784 5448 17584 5568
rect 0 2728 800 2848
rect 16784 2456 17584 2576
<< obsm3 >>
rect 800 17344 16784 17441
rect 880 17072 16784 17344
rect 880 17064 16704 17072
rect 800 16792 16704 17064
rect 800 14352 16784 16792
rect 880 14080 16784 14352
rect 880 14072 16704 14080
rect 800 13800 16704 14072
rect 800 11632 16784 13800
rect 880 11360 16784 11632
rect 880 11352 16704 11360
rect 800 11080 16704 11352
rect 800 8640 16784 11080
rect 880 8368 16784 8640
rect 880 8360 16704 8368
rect 800 8088 16704 8360
rect 800 5920 16784 8088
rect 880 5648 16784 5920
rect 880 5640 16704 5648
rect 800 5368 16704 5640
rect 800 2928 16784 5368
rect 880 2656 16784 2928
rect 880 2648 16704 2656
rect 800 2376 16704 2648
rect 800 2143 16784 2376
<< obsm4 >>
rect 3504 2128 14067 17456
<< metal5 >>
rect 1104 7046 16468 7366
rect 1104 4506 16468 4826
<< obsm5 >>
rect 1104 7686 16468 14981
<< labels >>
rlabel metal2 s 17498 18928 17554 19728 6 A[0]
port 1 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 A[1]
port 2 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 A[2]
port 3 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 A[3]
port 4 nsew signal input
rlabel metal2 s 5906 18928 5962 19728 6 A[4]
port 5 nsew signal input
rlabel metal2 s 11794 18928 11850 19728 6 A[5]
port 6 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 A[6]
port 7 nsew signal input
rlabel metal3 s 16784 8168 17584 8288 6 A[7]
port 8 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 B[0]
port 9 nsew signal input
rlabel metal3 s 16784 11160 17584 11280 6 B[1]
port 10 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 B[2]
port 11 nsew signal input
rlabel metal2 s 18 0 74 800 6 B[3]
port 12 nsew signal input
rlabel metal2 s 13634 18928 13690 19728 6 B[4]
port 13 nsew signal input
rlabel metal2 s 15658 18928 15714 19728 6 B[5]
port 14 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 B[6]
port 15 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 B[7]
port 16 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 M[0]
port 17 nsew signal output
rlabel metal2 s 18 18928 74 19728 6 M[10]
port 18 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 M[11]
port 19 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 M[12]
port 20 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 M[13]
port 21 nsew signal output
rlabel metal2 s 4066 18928 4122 19728 6 M[14]
port 22 nsew signal output
rlabel metal3 s 16784 2456 17584 2576 6 M[15]
port 23 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 M[1]
port 24 nsew signal output
rlabel metal3 s 16784 13880 17584 14000 6 M[2]
port 25 nsew signal output
rlabel metal3 s 16784 16872 17584 16992 6 M[3]
port 26 nsew signal output
rlabel metal2 s 7930 18928 7986 19728 6 M[4]
port 27 nsew signal output
rlabel metal2 s 9770 18928 9826 19728 6 M[5]
port 28 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 M[6]
port 29 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 M[7]
port 30 nsew signal output
rlabel metal2 s 2042 18928 2098 19728 6 M[8]
port 31 nsew signal output
rlabel metal3 s 16784 5448 17584 5568 6 M[9]
port 32 nsew signal output
rlabel metal5 s 1104 7046 16468 7366 6 VGND
port 33 nsew ground input
rlabel metal5 s 1104 4506 16468 4826 6 VPWR
port 34 nsew power input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 17584 19728
string LEFview TRUE
string GDS_FILE /openLANE_flow/designs/dvsd_8216m9/runs/20-08_18-30/results/magic/dvsd_8216m9.gds
string GDS_END 1167544
string GDS_START 224772
<< end >>


magic
tech sky130A
magscale 1 2
timestamp 1629722742
<< checkpaint >>
rect -3932 -3932 20803 22947
<< locali >>
rect 8769 10047 8803 10149
rect 5457 9911 5491 10013
rect 5825 8891 5859 9129
rect 10885 8959 10919 9129
rect 5549 6103 5583 6205
rect 10517 6171 10551 6341
<< viali >>
rect 4905 16133 4939 16167
rect 7665 16133 7699 16167
rect 9965 16133 9999 16167
rect 13277 16133 13311 16167
rect 1409 16065 1443 16099
rect 2881 16065 2915 16099
rect 2973 16065 3007 16099
rect 3249 16065 3283 16099
rect 4353 16065 4387 16099
rect 5089 16065 5123 16099
rect 6377 16065 6411 16099
rect 7849 16065 7883 16099
rect 9137 16065 9171 16099
rect 9229 16065 9263 16099
rect 9505 16065 9539 16099
rect 10149 16065 10183 16099
rect 11529 16065 11563 16099
rect 12541 16065 12575 16099
rect 14289 16065 14323 16099
rect 14841 16065 14875 16099
rect 15025 16065 15059 16099
rect 1685 15997 1719 16031
rect 6653 15997 6687 16031
rect 4169 15929 4203 15963
rect 12725 15929 12759 15963
rect 2697 15861 2731 15895
rect 3157 15861 3191 15895
rect 8953 15861 8987 15895
rect 9413 15861 9447 15895
rect 11713 15861 11747 15895
rect 13369 15861 13403 15895
rect 14105 15861 14139 15895
rect 9413 15657 9447 15691
rect 14657 15657 14691 15691
rect 8125 15589 8159 15623
rect 11161 15589 11195 15623
rect 12909 15589 12943 15623
rect 1501 15521 1535 15555
rect 2053 15521 2087 15555
rect 2697 15521 2731 15555
rect 3249 15521 3283 15555
rect 4537 15521 4571 15555
rect 4997 15521 5031 15555
rect 5733 15521 5767 15555
rect 9965 15521 9999 15555
rect 14933 15521 14967 15555
rect 1685 15453 1719 15487
rect 2881 15453 2915 15487
rect 4721 15453 4755 15487
rect 4813 15453 4847 15487
rect 5089 15453 5123 15487
rect 5825 15453 5859 15487
rect 7573 15453 7607 15487
rect 7849 15453 7883 15487
rect 7941 15453 7975 15487
rect 9597 15453 9631 15487
rect 9689 15453 9723 15487
rect 10609 15453 10643 15487
rect 10885 15453 10919 15487
rect 10977 15453 11011 15487
rect 11621 15453 11655 15487
rect 12357 15453 12391 15487
rect 12633 15453 12667 15487
rect 12725 15453 12759 15487
rect 13369 15453 13403 15487
rect 13553 15453 13587 15487
rect 14381 15453 14415 15487
rect 14749 15453 14783 15487
rect 1961 15385 1995 15419
rect 6101 15385 6135 15419
rect 6193 15385 6227 15419
rect 7481 15385 7515 15419
rect 10057 15385 10091 15419
rect 10517 15385 10551 15419
rect 12265 15385 12299 15419
rect 14473 15385 14507 15419
rect 1869 15317 1903 15351
rect 3065 15317 3099 15351
rect 3157 15317 3191 15351
rect 5549 15317 5583 15351
rect 11805 15317 11839 15351
rect 13461 15317 13495 15351
rect 2513 15113 2547 15147
rect 3433 15113 3467 15147
rect 5365 15113 5399 15147
rect 7113 15113 7147 15147
rect 9321 15113 9355 15147
rect 9413 15113 9447 15147
rect 12909 15113 12943 15147
rect 14473 15113 14507 15147
rect 2605 15045 2639 15079
rect 12817 15045 12851 15079
rect 1593 14977 1627 15011
rect 1685 14977 1719 15011
rect 1961 14977 1995 15011
rect 3709 14977 3743 15011
rect 3985 14977 4019 15011
rect 5641 14977 5675 15011
rect 7297 14977 7331 15011
rect 7389 14977 7423 15011
rect 7665 14977 7699 15011
rect 9597 14977 9631 15011
rect 9781 14977 9815 15011
rect 11621 14977 11655 15011
rect 11805 14977 11839 15011
rect 11897 14977 11931 15011
rect 12173 14977 12207 15011
rect 13093 14977 13127 15011
rect 14197 14977 14231 15011
rect 3617 14909 3651 14943
rect 4077 14909 4111 14943
rect 5273 14909 5307 14943
rect 5825 14909 5859 14943
rect 9229 14909 9263 14943
rect 12081 14909 12115 14943
rect 12725 14909 12759 14943
rect 13277 14909 13311 14943
rect 13829 14909 13863 14943
rect 13921 14909 13955 14943
rect 14289 14909 14323 14943
rect 1409 14773 1443 14807
rect 1869 14773 1903 14807
rect 5549 14773 5583 14807
rect 7573 14773 7607 14807
rect 1685 14569 1719 14603
rect 4537 14569 4571 14603
rect 7021 14569 7055 14603
rect 8953 14569 8987 14603
rect 10425 14569 10459 14603
rect 13001 14569 13035 14603
rect 14105 14569 14139 14603
rect 4997 14501 5031 14535
rect 12541 14501 12575 14535
rect 14565 14501 14599 14535
rect 1869 14433 1903 14467
rect 7205 14433 7239 14467
rect 10609 14433 10643 14467
rect 1961 14365 1995 14399
rect 4721 14365 4755 14399
rect 4813 14365 4847 14399
rect 5089 14365 5123 14399
rect 7297 14365 7331 14399
rect 7665 14365 7699 14399
rect 8309 14365 8343 14399
rect 9965 14365 9999 14399
rect 10701 14365 10735 14399
rect 11805 14365 11839 14399
rect 12449 14365 12483 14399
rect 12725 14365 12759 14399
rect 12817 14365 12851 14399
rect 14289 14365 14323 14399
rect 14381 14365 14415 14399
rect 14657 14365 14691 14399
rect 2237 14297 2271 14331
rect 2329 14297 2363 14331
rect 7573 14297 7607 14331
rect 9137 14297 9171 14331
rect 9321 14297 9355 14331
rect 10977 14297 11011 14331
rect 11069 14297 11103 14331
rect 8217 14229 8251 14263
rect 9781 14229 9815 14263
rect 11897 14229 11931 14263
rect 3157 14025 3191 14059
rect 4813 14025 4847 14059
rect 7849 14025 7883 14059
rect 10333 14025 10367 14059
rect 13461 14025 13495 14059
rect 2053 13957 2087 13991
rect 9689 13957 9723 13991
rect 1869 13889 1903 13923
rect 2605 13889 2639 13923
rect 2881 13889 2915 13923
rect 5089 13889 5123 13923
rect 5365 13889 5399 13923
rect 6929 13889 6963 13923
rect 8125 13889 8159 13923
rect 8401 13889 8435 13923
rect 9505 13889 9539 13923
rect 9873 13889 9907 13923
rect 10517 13889 10551 13923
rect 10609 13889 10643 13923
rect 10885 13889 10919 13923
rect 11713 13889 11747 13923
rect 12173 13889 12207 13923
rect 12817 13889 12851 13923
rect 13185 13889 13219 13923
rect 14105 13889 14139 13923
rect 14841 13889 14875 13923
rect 2513 13821 2547 13855
rect 2973 13821 3007 13855
rect 4997 13821 5031 13855
rect 5457 13821 5491 13855
rect 8033 13821 8067 13855
rect 8493 13821 8527 13855
rect 10793 13821 10827 13855
rect 12909 13821 12943 13855
rect 13277 13821 13311 13855
rect 14197 13821 14231 13855
rect 15025 13821 15059 13855
rect 7113 13685 7147 13719
rect 11621 13685 11655 13719
rect 12357 13685 12391 13719
rect 2697 13481 2731 13515
rect 5549 13481 5583 13515
rect 7205 13481 7239 13515
rect 7389 13481 7423 13515
rect 8953 13481 8987 13515
rect 11161 13481 11195 13515
rect 12541 13481 12575 13515
rect 13369 13481 13403 13515
rect 14749 13481 14783 13515
rect 7849 13413 7883 13447
rect 14289 13413 14323 13447
rect 2237 13345 2271 13379
rect 4997 13345 5031 13379
rect 8309 13345 8343 13379
rect 9597 13345 9631 13379
rect 11989 13345 12023 13379
rect 12357 13345 12391 13379
rect 2145 13277 2179 13311
rect 2421 13277 2455 13311
rect 2513 13277 2547 13311
rect 5273 13277 5307 13311
rect 5365 13277 5399 13311
rect 6929 13277 6963 13311
rect 8033 13277 8067 13311
rect 8125 13277 8159 13311
rect 8401 13277 8435 13311
rect 9137 13277 9171 13311
rect 9229 13277 9263 13311
rect 9505 13277 9539 13311
rect 10517 13277 10551 13311
rect 11191 13277 11225 13311
rect 11345 13277 11379 13311
rect 12265 13277 12299 13311
rect 13185 13277 13219 13311
rect 14197 13277 14231 13311
rect 14473 13277 14507 13311
rect 14565 13277 14599 13311
rect 4905 13209 4939 13243
rect 11897 13209 11931 13243
rect 13001 13209 13035 13243
rect 10333 13141 10367 13175
rect 2237 12937 2271 12971
rect 3525 12937 3559 12971
rect 5733 12937 5767 12971
rect 11989 12937 12023 12971
rect 14749 12937 14783 12971
rect 1593 12869 1627 12903
rect 2973 12869 3007 12903
rect 1961 12801 1995 12835
rect 2881 12801 2915 12835
rect 3249 12801 3283 12835
rect 4261 12801 4295 12835
rect 5825 12801 5859 12835
rect 6561 12801 6595 12835
rect 7481 12801 7515 12835
rect 9229 12801 9263 12835
rect 9413 12801 9447 12835
rect 9965 12801 9999 12835
rect 10241 12801 10275 12835
rect 10333 12801 10367 12835
rect 11529 12801 11563 12835
rect 11805 12801 11839 12835
rect 12449 12801 12483 12835
rect 13185 12801 13219 12835
rect 14473 12801 14507 12835
rect 1685 12733 1719 12767
rect 2053 12733 2087 12767
rect 3341 12733 3375 12767
rect 4169 12733 4203 12767
rect 4537 12733 4571 12767
rect 4629 12733 4663 12767
rect 7757 12733 7791 12767
rect 11621 12733 11655 12767
rect 13645 12733 13679 12767
rect 14105 12733 14139 12767
rect 14197 12733 14231 12767
rect 14565 12733 14599 12767
rect 10517 12665 10551 12699
rect 3985 12597 4019 12631
rect 6653 12597 6687 12631
rect 9045 12597 9079 12631
rect 10057 12597 10091 12631
rect 11805 12597 11839 12631
rect 12633 12597 12667 12631
rect 13277 12597 13311 12631
rect 3801 12393 3835 12427
rect 5365 12393 5399 12427
rect 7205 12393 7239 12427
rect 7665 12393 7699 12427
rect 8217 12393 8251 12427
rect 9229 12393 9263 12427
rect 10241 12393 10275 12427
rect 11897 12393 11931 12427
rect 13553 12393 13587 12427
rect 14749 12393 14783 12427
rect 10701 12325 10735 12359
rect 4261 12257 4295 12291
rect 9689 12257 9723 12291
rect 10333 12257 10367 12291
rect 14473 12257 14507 12291
rect 15025 12257 15059 12291
rect 3985 12189 4019 12223
rect 4077 12189 4111 12223
rect 4353 12189 4387 12223
rect 5549 12189 5583 12223
rect 5641 12189 5675 12223
rect 5917 12189 5951 12223
rect 6561 12189 6595 12223
rect 7389 12189 7423 12223
rect 7481 12189 7515 12223
rect 7757 12189 7791 12223
rect 8401 12189 8435 12223
rect 9413 12189 9447 12223
rect 9505 12189 9539 12223
rect 9781 12189 9815 12223
rect 10517 12189 10551 12223
rect 11713 12189 11747 12223
rect 13185 12189 13219 12223
rect 13369 12189 13403 12223
rect 14841 12189 14875 12223
rect 6009 12121 6043 12155
rect 10241 12121 10275 12155
rect 11529 12121 11563 12155
rect 12357 12121 12391 12155
rect 12541 12121 12575 12155
rect 6745 12053 6779 12087
rect 12725 12053 12759 12087
rect 14565 12053 14599 12087
rect 1685 11849 1719 11883
rect 7205 11849 7239 11883
rect 8033 11849 8067 11883
rect 10149 11849 10183 11883
rect 10793 11849 10827 11883
rect 11529 11849 11563 11883
rect 4353 11781 4387 11815
rect 6745 11781 6779 11815
rect 8861 11781 8895 11815
rect 12909 11781 12943 11815
rect 1961 11713 1995 11747
rect 2237 11713 2271 11747
rect 3617 11713 3651 11747
rect 3801 11713 3835 11747
rect 3893 11713 3927 11747
rect 4537 11713 4571 11747
rect 4721 11713 4755 11747
rect 5365 11713 5399 11747
rect 5594 11713 5628 11747
rect 5825 11713 5859 11747
rect 7021 11713 7055 11747
rect 7849 11713 7883 11747
rect 8493 11713 8527 11747
rect 8677 11713 8711 11747
rect 9321 11713 9355 11747
rect 9505 11713 9539 11747
rect 10333 11713 10367 11747
rect 10977 11713 11011 11747
rect 11713 11713 11747 11747
rect 11805 11713 11839 11747
rect 12081 11713 12115 11747
rect 13185 11713 13219 11747
rect 14105 11713 14139 11747
rect 14933 11713 14967 11747
rect 1869 11645 1903 11679
rect 2329 11645 2363 11679
rect 6837 11645 6871 11679
rect 12817 11645 12851 11679
rect 13277 11645 13311 11679
rect 14197 11645 14231 11679
rect 5181 11577 5215 11611
rect 14749 11577 14783 11611
rect 3617 11509 3651 11543
rect 6837 11509 6871 11543
rect 9321 11509 9355 11543
rect 11989 11509 12023 11543
rect 13461 11509 13495 11543
rect 1501 11305 1535 11339
rect 2697 11305 2731 11339
rect 3801 11305 3835 11339
rect 5273 11305 5307 11339
rect 6561 11305 6595 11339
rect 10977 11305 11011 11339
rect 11161 11305 11195 11339
rect 12725 11305 12759 11339
rect 13185 11305 13219 11339
rect 14105 11305 14139 11339
rect 5825 11237 5859 11271
rect 7021 11237 7055 11271
rect 10241 11237 10275 11271
rect 12265 11237 12299 11271
rect 1685 11169 1719 11203
rect 2145 11169 2179 11203
rect 4445 11169 4479 11203
rect 7573 11169 7607 11203
rect 11345 11169 11379 11203
rect 14289 11169 14323 11203
rect 14749 11169 14783 11203
rect 1777 11101 1811 11135
rect 2605 11101 2639 11135
rect 2821 11101 2855 11135
rect 2973 11101 3007 11135
rect 3985 11101 4019 11135
rect 4077 11101 4111 11135
rect 5641 11101 5675 11135
rect 6745 11101 6779 11135
rect 6837 11101 6871 11135
rect 7113 11101 7147 11135
rect 7849 11101 7883 11135
rect 9137 11101 9171 11135
rect 11161 11101 11195 11135
rect 11897 11101 11931 11135
rect 12051 11101 12085 11135
rect 12909 11101 12943 11135
rect 13001 11101 13035 11135
rect 13277 11101 13311 11135
rect 14381 11101 14415 11135
rect 14657 11101 14691 11135
rect 2053 11033 2087 11067
rect 3157 11033 3191 11067
rect 4353 11033 4387 11067
rect 5549 11033 5583 11067
rect 9873 11033 9907 11067
rect 10057 11033 10091 11067
rect 11437 11033 11471 11067
rect 5457 10965 5491 10999
rect 8953 10965 8987 10999
rect 2053 10761 2087 10795
rect 3617 10761 3651 10795
rect 4353 10761 4387 10795
rect 6469 10761 6503 10795
rect 9229 10761 9263 10795
rect 4169 10693 4203 10727
rect 4445 10693 4479 10727
rect 5457 10693 5491 10727
rect 9781 10693 9815 10727
rect 10517 10693 10551 10727
rect 13921 10693 13955 10727
rect 14565 10693 14599 10727
rect 2237 10625 2271 10659
rect 2329 10625 2363 10659
rect 2605 10625 2639 10659
rect 3525 10625 3559 10659
rect 3709 10625 3743 10659
rect 4537 10625 4571 10659
rect 5641 10625 5675 10659
rect 6377 10625 6411 10659
rect 6561 10625 6595 10659
rect 7205 10625 7239 10659
rect 7297 10625 7331 10659
rect 7573 10625 7607 10659
rect 8033 10625 8067 10659
rect 8309 10625 8343 10659
rect 9505 10625 9539 10659
rect 10701 10625 10735 10659
rect 11713 10625 11747 10659
rect 12449 10625 12483 10659
rect 12541 10625 12575 10659
rect 13001 10625 13035 10659
rect 13185 10625 13219 10659
rect 13737 10625 13771 10659
rect 7021 10557 7055 10591
rect 7481 10557 7515 10591
rect 8125 10557 8159 10591
rect 9413 10557 9447 10591
rect 9873 10557 9907 10591
rect 10333 10557 10367 10591
rect 14381 10557 14415 10591
rect 4721 10489 4755 10523
rect 5825 10489 5859 10523
rect 13185 10489 13219 10523
rect 2513 10421 2547 10455
rect 8125 10421 8159 10455
rect 8493 10421 8527 10455
rect 11529 10421 11563 10455
rect 1869 10217 1903 10251
rect 3157 10217 3191 10251
rect 4077 10217 4111 10251
rect 7849 10217 7883 10251
rect 10793 10217 10827 10251
rect 11989 10217 12023 10251
rect 13185 10217 13219 10251
rect 8769 10149 8803 10183
rect 11253 10149 11287 10183
rect 12449 10149 12483 10183
rect 4629 10081 4663 10115
rect 14105 10081 14139 10115
rect 1961 10013 1995 10047
rect 2881 10013 2915 10047
rect 2973 10013 3007 10047
rect 4169 10013 4203 10047
rect 4873 10013 4907 10047
rect 4997 10013 5031 10047
rect 5457 10013 5491 10047
rect 5549 10013 5583 10047
rect 6653 10013 6687 10047
rect 7849 10013 7883 10047
rect 7941 10013 7975 10047
rect 8125 10013 8159 10047
rect 8769 10013 8803 10047
rect 9137 10013 9171 10047
rect 9321 10013 9355 10047
rect 9597 10013 9631 10047
rect 9781 10013 9815 10047
rect 10977 10013 11011 10047
rect 11069 10013 11103 10047
rect 11345 10013 11379 10047
rect 12173 10013 12207 10047
rect 12265 10013 12299 10047
rect 12541 10013 12575 10047
rect 13185 10013 13219 10047
rect 13277 10013 13311 10047
rect 14381 10013 14415 10047
rect 2513 9945 2547 9979
rect 2605 9945 2639 9979
rect 6285 9945 6319 9979
rect 6469 9945 6503 9979
rect 13001 9945 13035 9979
rect 5457 9877 5491 9911
rect 5641 9877 5675 9911
rect 7665 9877 7699 9911
rect 13461 9877 13495 9911
rect 2053 9673 2087 9707
rect 9505 9673 9539 9707
rect 9873 9673 9907 9707
rect 10609 9673 10643 9707
rect 11621 9673 11655 9707
rect 9689 9605 9723 9639
rect 12081 9605 12115 9639
rect 2329 9537 2363 9571
rect 2605 9537 2639 9571
rect 3985 9537 4019 9571
rect 4077 9537 4111 9571
rect 5089 9537 5123 9571
rect 5181 9537 5215 9571
rect 5549 9537 5583 9571
rect 6838 9537 6872 9571
rect 6989 9537 7023 9571
rect 7205 9537 7239 9571
rect 7757 9537 7791 9571
rect 9781 9537 9815 9571
rect 10517 9537 10551 9571
rect 11805 9537 11839 9571
rect 13277 9537 13311 9571
rect 14657 9537 14691 9571
rect 14749 9537 14783 9571
rect 2237 9469 2271 9503
rect 2697 9469 2731 9503
rect 4353 9469 4387 9503
rect 4445 9469 4479 9503
rect 5457 9469 5491 9503
rect 8033 9469 8067 9503
rect 11897 9469 11931 9503
rect 12909 9469 12943 9503
rect 14381 9469 14415 9503
rect 14565 9469 14599 9503
rect 14841 9469 14875 9503
rect 3801 9401 3835 9435
rect 4905 9401 4939 9435
rect 10057 9401 10091 9435
rect 6653 9333 6687 9367
rect 7113 9333 7147 9367
rect 11805 9333 11839 9367
rect 2329 9129 2363 9163
rect 4905 9129 4939 9163
rect 5825 9129 5859 9163
rect 6009 9129 6043 9163
rect 6377 9129 6411 9163
rect 7849 9129 7883 9163
rect 9321 9129 9355 9163
rect 10885 9129 10919 9163
rect 12817 9129 12851 9163
rect 14473 9129 14507 9163
rect 3249 9061 3283 9095
rect 1685 8993 1719 9027
rect 2053 8925 2087 8959
rect 2145 8925 2179 8959
rect 3065 8925 3099 8959
rect 3801 8925 3835 8959
rect 4629 8925 4663 8959
rect 4721 8925 4755 8959
rect 4997 8925 5031 8959
rect 6469 8925 6503 8959
rect 7573 8925 7607 8959
rect 7665 8925 7699 8959
rect 7941 8925 7975 8959
rect 9781 8925 9815 8959
rect 9965 8925 9999 8959
rect 10885 8925 10919 8959
rect 11161 8925 11195 8959
rect 11621 8925 11655 8959
rect 13093 8925 13127 8959
rect 14105 8925 14139 8959
rect 14289 8925 14323 8959
rect 1777 8857 1811 8891
rect 5825 8857 5859 8891
rect 8953 8857 8987 8891
rect 9137 8857 9171 8891
rect 11805 8857 11839 8891
rect 3985 8789 4019 8823
rect 4445 8789 4479 8823
rect 7389 8789 7423 8823
rect 9873 8789 9907 8823
rect 11069 8789 11103 8823
rect 11989 8789 12023 8823
rect 9321 8585 9355 8619
rect 11529 8585 11563 8619
rect 14565 8585 14599 8619
rect 4261 8517 4295 8551
rect 5825 8517 5859 8551
rect 9873 8517 9907 8551
rect 14749 8517 14783 8551
rect 1961 8449 1995 8483
rect 2053 8449 2087 8483
rect 2421 8449 2455 8483
rect 3065 8449 3099 8483
rect 3801 8449 3835 8483
rect 3893 8449 3927 8483
rect 4169 8449 4203 8483
rect 5365 8449 5399 8483
rect 5457 8449 5491 8483
rect 6469 8449 6503 8483
rect 7573 8449 7607 8483
rect 8861 8449 8895 8483
rect 9597 8449 9631 8483
rect 10425 8449 10459 8483
rect 10609 8449 10643 8483
rect 11713 8449 11747 8483
rect 11805 8449 11839 8483
rect 12081 8449 12115 8483
rect 13093 8449 13127 8483
rect 13277 8449 13311 8483
rect 13737 8449 13771 8483
rect 13829 8449 13863 8483
rect 14473 8449 14507 8483
rect 2329 8381 2363 8415
rect 5733 8381 5767 8415
rect 8585 8381 8619 8415
rect 9505 8381 9539 8415
rect 9965 8381 9999 8415
rect 10517 8381 10551 8415
rect 14013 8381 14047 8415
rect 2881 8313 2915 8347
rect 7113 8313 7147 8347
rect 11989 8313 12023 8347
rect 13921 8313 13955 8347
rect 14749 8313 14783 8347
rect 1777 8245 1811 8279
rect 3617 8245 3651 8279
rect 5181 8245 5215 8279
rect 6561 8245 6595 8279
rect 7389 8245 7423 8279
rect 12909 8245 12943 8279
rect 2053 8041 2087 8075
rect 2605 8041 2639 8075
rect 3985 8041 4019 8075
rect 10885 8041 10919 8075
rect 12633 8041 12667 8075
rect 4445 7973 4479 8007
rect 9321 7973 9355 8007
rect 13185 7973 13219 8007
rect 2789 7905 2823 7939
rect 3157 7905 3191 7939
rect 3249 7905 3283 7939
rect 4997 7905 5031 7939
rect 11345 7905 11379 7939
rect 1777 7837 1811 7871
rect 1869 7837 1903 7871
rect 2145 7837 2179 7871
rect 2881 7837 2915 7871
rect 3801 7837 3835 7871
rect 3985 7837 4019 7871
rect 4629 7837 4663 7871
rect 4721 7837 4755 7871
rect 6286 7847 6320 7881
rect 6745 7837 6779 7871
rect 7205 7837 7239 7871
rect 8401 7837 8435 7871
rect 9321 7837 9355 7871
rect 9597 7837 9631 7871
rect 10425 7837 10459 7871
rect 11069 7837 11103 7871
rect 11161 7837 11195 7871
rect 11437 7837 11471 7871
rect 11989 7837 12023 7871
rect 12909 7837 12943 7871
rect 14197 7837 14231 7871
rect 14473 7837 14507 7871
rect 5089 7769 5123 7803
rect 6377 7769 6411 7803
rect 6469 7769 6503 7803
rect 6607 7769 6641 7803
rect 7297 7769 7331 7803
rect 9505 7769 9539 7803
rect 12817 7769 12851 7803
rect 1593 7701 1627 7735
rect 6101 7701 6135 7735
rect 8217 7701 8251 7735
rect 10333 7701 10367 7735
rect 12173 7701 12207 7735
rect 13001 7701 13035 7735
rect 2973 7497 3007 7531
rect 6929 7497 6963 7531
rect 13461 7497 13495 7531
rect 12541 7429 12575 7463
rect 12771 7429 12805 7463
rect 2881 7361 2915 7395
rect 3709 7361 3743 7395
rect 3801 7361 3835 7395
rect 4077 7361 4111 7395
rect 5273 7361 5307 7395
rect 5365 7361 5399 7395
rect 5641 7361 5675 7395
rect 7113 7361 7147 7395
rect 7389 7361 7423 7395
rect 7573 7361 7607 7395
rect 8217 7361 8251 7395
rect 9137 7361 9171 7395
rect 9781 7361 9815 7395
rect 10333 7361 10367 7395
rect 11621 7361 11655 7395
rect 12449 7361 12483 7395
rect 12633 7361 12667 7395
rect 13369 7361 13403 7395
rect 14197 7361 14231 7395
rect 14473 7361 14507 7395
rect 3985 7293 4019 7327
rect 7297 7293 7331 7327
rect 12909 7293 12943 7327
rect 14289 7293 14323 7327
rect 14381 7293 14415 7327
rect 7205 7225 7239 7259
rect 8125 7225 8159 7259
rect 9045 7225 9079 7259
rect 3525 7157 3559 7191
rect 5089 7157 5123 7191
rect 5549 7157 5583 7191
rect 9597 7157 9631 7191
rect 10425 7157 10459 7191
rect 11805 7157 11839 7191
rect 12265 7157 12299 7191
rect 14013 7157 14047 7191
rect 10977 6953 11011 6987
rect 13185 6953 13219 6987
rect 12541 6885 12575 6919
rect 4261 6817 4295 6851
rect 5089 6817 5123 6851
rect 5549 6817 5583 6851
rect 6193 6817 6227 6851
rect 6561 6817 6595 6851
rect 7665 6817 7699 6851
rect 8309 6817 8343 6851
rect 11529 6817 11563 6851
rect 14105 6817 14139 6851
rect 14381 6817 14415 6851
rect 1869 6749 1903 6783
rect 2053 6749 2087 6783
rect 2421 6749 2455 6783
rect 3985 6749 4019 6783
rect 4077 6749 4111 6783
rect 4353 6749 4387 6783
rect 5181 6749 5215 6783
rect 5457 6749 5491 6783
rect 6377 6749 6411 6783
rect 6469 6749 6503 6783
rect 6653 6749 6687 6783
rect 6837 6749 6871 6783
rect 7573 6749 7607 6783
rect 7757 6749 7791 6783
rect 8217 6749 8251 6783
rect 8401 6749 8435 6783
rect 9137 6749 9171 6783
rect 9229 6749 9263 6783
rect 9505 6749 9539 6783
rect 10149 6749 10183 6783
rect 11130 6749 11164 6783
rect 11621 6749 11655 6783
rect 12265 6749 12299 6783
rect 12357 6749 12391 6783
rect 12633 6749 12667 6783
rect 13093 6749 13127 6783
rect 9597 6681 9631 6715
rect 10333 6681 10367 6715
rect 10517 6681 10551 6715
rect 11226 6681 11260 6715
rect 2145 6613 2179 6647
rect 2329 6613 2363 6647
rect 3801 6613 3835 6647
rect 4905 6613 4939 6647
rect 8953 6613 8987 6647
rect 12081 6613 12115 6647
rect 1869 6409 1903 6443
rect 3985 6409 4019 6443
rect 4445 6409 4479 6443
rect 7941 6409 7975 6443
rect 9597 6409 9631 6443
rect 3341 6341 3375 6375
rect 5089 6341 5123 6375
rect 7021 6341 7055 6375
rect 7113 6341 7147 6375
rect 8493 6341 8527 6375
rect 9689 6341 9723 6375
rect 10517 6341 10551 6375
rect 10609 6341 10643 6375
rect 2145 6273 2179 6307
rect 3433 6273 3467 6307
rect 3709 6273 3743 6307
rect 4629 6273 4663 6307
rect 4721 6273 4755 6307
rect 5641 6273 5675 6307
rect 5825 6273 5859 6307
rect 6929 6273 6963 6307
rect 8217 6273 8251 6307
rect 9505 6273 9539 6307
rect 1777 6205 1811 6239
rect 2329 6205 2363 6239
rect 3801 6205 3835 6239
rect 4997 6205 5031 6239
rect 5549 6205 5583 6239
rect 8125 6205 8159 6239
rect 8585 6205 8619 6239
rect 10793 6273 10827 6307
rect 11805 6273 11839 6307
rect 11989 6273 12023 6307
rect 12817 6273 12851 6307
rect 12909 6273 12943 6307
rect 13001 6273 13035 6307
rect 13139 6273 13173 6307
rect 13829 6273 13863 6307
rect 14105 6273 14139 6307
rect 14289 6273 14323 6307
rect 11713 6205 11747 6239
rect 13277 6205 13311 6239
rect 14013 6205 14047 6239
rect 14197 6205 14231 6239
rect 7297 6137 7331 6171
rect 9321 6137 9355 6171
rect 9873 6137 9907 6171
rect 10517 6137 10551 6171
rect 2053 6069 2087 6103
rect 5549 6069 5583 6103
rect 5641 6069 5675 6103
rect 6745 6069 6779 6103
rect 10977 6069 11011 6103
rect 12173 6069 12207 6103
rect 12633 6069 12667 6103
rect 14473 6069 14507 6103
rect 8309 5865 8343 5899
rect 11529 5865 11563 5899
rect 13461 5865 13495 5899
rect 14841 5865 14875 5899
rect 3249 5797 3283 5831
rect 5733 5797 5767 5831
rect 7113 5797 7147 5831
rect 9505 5797 9539 5831
rect 10057 5797 10091 5831
rect 10977 5797 11011 5831
rect 1869 5729 1903 5763
rect 3985 5729 4019 5763
rect 4445 5729 4479 5763
rect 5917 5729 5951 5763
rect 6377 5729 6411 5763
rect 9321 5729 9355 5763
rect 14381 5729 14415 5763
rect 14473 5729 14507 5763
rect 1593 5661 1627 5695
rect 1685 5661 1719 5695
rect 1961 5661 1995 5695
rect 2421 5661 2455 5695
rect 3065 5661 3099 5695
rect 4077 5661 4111 5695
rect 4353 5661 4387 5695
rect 5273 5661 5307 5695
rect 6009 5661 6043 5695
rect 6285 5661 6319 5695
rect 6837 5661 6871 5695
rect 6929 5661 6963 5695
rect 8033 5661 8067 5695
rect 8125 5661 8159 5695
rect 8401 5661 8435 5695
rect 9597 5661 9631 5695
rect 10342 5661 10376 5695
rect 10793 5661 10827 5695
rect 10977 5661 11011 5695
rect 11437 5661 11471 5695
rect 11621 5661 11655 5695
rect 12081 5661 12115 5695
rect 12265 5661 12299 5695
rect 12909 5661 12943 5695
rect 13553 5661 13587 5695
rect 14657 5661 14691 5695
rect 7113 5593 7147 5627
rect 9321 5593 9355 5627
rect 10057 5593 10091 5627
rect 1409 5525 1443 5559
rect 2605 5525 2639 5559
rect 3801 5525 3835 5559
rect 5181 5525 5215 5559
rect 7849 5525 7883 5559
rect 10241 5525 10275 5559
rect 12173 5525 12207 5559
rect 12817 5525 12851 5559
rect 1593 5321 1627 5355
rect 2605 5321 2639 5355
rect 7021 5321 7055 5355
rect 10517 5321 10551 5355
rect 11621 5321 11655 5355
rect 13185 5321 13219 5355
rect 14197 5321 14231 5355
rect 14841 5253 14875 5287
rect 1409 5185 1443 5219
rect 2421 5185 2455 5219
rect 3065 5185 3099 5219
rect 3893 5185 3927 5219
rect 3985 5185 4019 5219
rect 4261 5185 4295 5219
rect 4721 5185 4755 5219
rect 4905 5185 4939 5219
rect 4997 5185 5031 5219
rect 5273 5185 5307 5219
rect 6929 5185 6963 5219
rect 7113 5185 7147 5219
rect 7757 5185 7791 5219
rect 7941 5185 7975 5219
rect 8033 5185 8067 5219
rect 8309 5185 8343 5219
rect 8769 5185 8803 5219
rect 9045 5185 9079 5219
rect 9137 5185 9171 5219
rect 10057 5185 10091 5219
rect 10149 5185 10183 5219
rect 10333 5185 10367 5219
rect 11805 5185 11839 5219
rect 11989 5185 12023 5219
rect 12081 5185 12115 5219
rect 12817 5185 12851 5219
rect 13001 5185 13035 5219
rect 14105 5185 14139 5219
rect 14289 5185 14323 5219
rect 15025 5185 15059 5219
rect 5181 5117 5215 5151
rect 10241 5117 10275 5151
rect 11897 5117 11931 5151
rect 3157 5049 3191 5083
rect 8861 5049 8895 5083
rect 3709 4981 3743 5015
rect 4169 4981 4203 5015
rect 8217 4981 8251 5015
rect 9321 4981 9355 5015
rect 1685 4777 1719 4811
rect 4169 4777 4203 4811
rect 8217 4777 8251 4811
rect 10241 4777 10275 4811
rect 2697 4709 2731 4743
rect 1409 4641 1443 4675
rect 1961 4641 1995 4675
rect 4353 4641 4387 4675
rect 4813 4641 4847 4675
rect 5825 4641 5859 4675
rect 6469 4641 6503 4675
rect 7297 4641 7331 4675
rect 7757 4641 7791 4675
rect 9413 4641 9447 4675
rect 9505 4641 9539 4675
rect 12909 4641 12943 4675
rect 14473 4641 14507 4675
rect 1593 4573 1627 4607
rect 2513 4573 2547 4607
rect 2605 4573 2639 4607
rect 3065 4573 3099 4607
rect 4445 4573 4479 4607
rect 4721 4573 4755 4607
rect 5457 4573 5491 4607
rect 5549 4573 5583 4607
rect 6377 4573 6411 4607
rect 6561 4573 6595 4607
rect 7389 4573 7423 4607
rect 7665 4573 7699 4607
rect 8401 4573 8435 4607
rect 9321 4573 9355 4607
rect 9600 4573 9634 4607
rect 10609 4573 10643 4607
rect 11437 4573 11471 4607
rect 11529 4573 11563 4607
rect 11897 4573 11931 4607
rect 13093 4573 13127 4607
rect 13277 4573 13311 4607
rect 13395 4573 13429 4607
rect 13553 4573 13587 4607
rect 14289 4573 14323 4607
rect 14565 4573 14599 4607
rect 14657 4573 14691 4607
rect 14749 4573 14783 4607
rect 1869 4505 1903 4539
rect 5917 4505 5951 4539
rect 10425 4505 10459 4539
rect 11621 4505 11655 4539
rect 11759 4505 11793 4539
rect 13185 4505 13219 4539
rect 2973 4437 3007 4471
rect 5273 4437 5307 4471
rect 7113 4437 7147 4471
rect 9781 4437 9815 4471
rect 11253 4437 11287 4471
rect 14933 4437 14967 4471
rect 3709 4233 3743 4267
rect 5181 4233 5215 4267
rect 6469 4233 6503 4267
rect 8953 4233 8987 4267
rect 14473 4233 14507 4267
rect 4353 4165 4387 4199
rect 11897 4165 11931 4199
rect 13093 4165 13127 4199
rect 2053 4097 2087 4131
rect 2145 4097 2179 4131
rect 2421 4097 2455 4131
rect 3249 4097 3283 4131
rect 3985 4097 4019 4131
rect 4261 4097 4295 4131
rect 5457 4097 5491 4131
rect 5733 4097 5767 4131
rect 6561 4097 6595 4131
rect 7021 4097 7055 4131
rect 7297 4097 7331 4131
rect 7389 4097 7423 4131
rect 8217 4097 8251 4131
rect 8401 4097 8435 4131
rect 8861 4097 8895 4131
rect 9045 4097 9079 4131
rect 9505 4097 9539 4131
rect 10149 4097 10183 4131
rect 10977 4097 11011 4131
rect 11713 4097 11747 4131
rect 11805 4097 11839 4131
rect 12081 4097 12115 4131
rect 12909 4097 12943 4131
rect 13829 4097 13863 4131
rect 14197 4097 14231 4131
rect 14289 4097 14323 4131
rect 2329 4029 2363 4063
rect 3893 4029 3927 4063
rect 5365 4029 5399 4063
rect 5825 4029 5859 4063
rect 10885 4029 10919 4063
rect 13277 4029 13311 4063
rect 14013 4029 14047 4063
rect 14105 4029 14139 4063
rect 7113 3961 7147 3995
rect 8401 3961 8435 3995
rect 11529 3961 11563 3995
rect 1869 3893 1903 3927
rect 3157 3893 3191 3927
rect 7573 3893 7607 3927
rect 9597 3893 9631 3927
rect 10241 3893 10275 3927
rect 14105 3689 14139 3723
rect 2145 3621 2179 3655
rect 5089 3621 5123 3655
rect 6377 3621 6411 3655
rect 9689 3621 9723 3655
rect 14381 3621 14415 3655
rect 1869 3553 1903 3587
rect 2421 3553 2455 3587
rect 4629 3553 4663 3587
rect 7113 3553 7147 3587
rect 9597 3553 9631 3587
rect 9965 3553 9999 3587
rect 11989 3553 12023 3587
rect 14473 3553 14507 3587
rect 14565 3553 14599 3587
rect 2053 3485 2087 3519
rect 3249 3485 3283 3519
rect 3985 3485 4019 3519
rect 4813 3485 4847 3519
rect 4905 3485 4939 3519
rect 5181 3485 5215 3519
rect 6193 3485 6227 3519
rect 7021 3485 7055 3519
rect 7205 3485 7239 3519
rect 7297 3485 7331 3519
rect 7481 3485 7515 3519
rect 7947 3485 7981 3519
rect 8125 3485 8159 3519
rect 9321 3485 9355 3519
rect 9505 3485 9539 3519
rect 9781 3485 9815 3519
rect 10885 3485 10919 3519
rect 11069 3485 11103 3519
rect 11253 3485 11287 3519
rect 11897 3485 11931 3519
rect 12173 3485 12207 3519
rect 12265 3485 12299 3519
rect 13369 3485 13403 3519
rect 14289 3485 14323 3519
rect 14749 3485 14783 3519
rect 3893 3417 3927 3451
rect 11161 3417 11195 3451
rect 13553 3417 13587 3451
rect 2329 3349 2363 3383
rect 3157 3349 3191 3383
rect 6837 3349 6871 3383
rect 8033 3349 8067 3383
rect 11437 3349 11471 3383
rect 12449 3349 12483 3383
rect 7757 3145 7791 3179
rect 8585 3145 8619 3179
rect 9229 3145 9263 3179
rect 9413 3145 9447 3179
rect 10333 3145 10367 3179
rect 11621 3145 11655 3179
rect 3801 3077 3835 3111
rect 5641 3077 5675 3111
rect 10885 3077 10919 3111
rect 2881 3009 2915 3043
rect 3617 3009 3651 3043
rect 3709 3009 3743 3043
rect 3985 3009 4019 3043
rect 4629 3009 4663 3043
rect 5457 3009 5491 3043
rect 5549 3009 5583 3043
rect 5825 3009 5859 3043
rect 6745 3009 6779 3043
rect 7297 3009 7331 3043
rect 7760 3009 7794 3043
rect 8677 3009 8711 3043
rect 9410 3009 9444 3043
rect 10609 3009 10643 3043
rect 11529 3009 11563 3043
rect 12173 3009 12207 3043
rect 12357 3009 12391 3043
rect 13001 3009 13035 3043
rect 13645 3009 13679 3043
rect 14013 3009 14047 3043
rect 14473 3009 14507 3043
rect 1409 2941 1443 2975
rect 1685 2941 1719 2975
rect 7389 2941 7423 2975
rect 9873 2941 9907 2975
rect 10517 2941 10551 2975
rect 10977 2941 11011 2975
rect 13093 2941 13127 2975
rect 14657 2941 14691 2975
rect 2697 2873 2731 2907
rect 4445 2873 4479 2907
rect 6561 2873 6595 2907
rect 12449 2873 12483 2907
rect 14197 2873 14231 2907
rect 3433 2805 3467 2839
rect 5273 2805 5307 2839
rect 7941 2805 7975 2839
rect 9781 2805 9815 2839
rect 3157 2601 3191 2635
rect 5089 2601 5123 2635
rect 8033 2601 8067 2635
rect 11621 2601 11655 2635
rect 13369 2601 13403 2635
rect 15025 2601 15059 2635
rect 4077 2533 4111 2567
rect 7113 2533 7147 2567
rect 12081 2533 12115 2567
rect 1685 2465 1719 2499
rect 3801 2465 3835 2499
rect 4353 2465 4387 2499
rect 4813 2465 4847 2499
rect 5365 2465 5399 2499
rect 7205 2465 7239 2499
rect 7297 2465 7331 2499
rect 9321 2465 9355 2499
rect 10885 2465 10919 2499
rect 12817 2465 12851 2499
rect 1409 2397 1443 2431
rect 2881 2397 2915 2431
rect 2973 2397 3007 2431
rect 3249 2397 3283 2431
rect 4169 2397 4203 2431
rect 5181 2397 5215 2431
rect 7021 2397 7055 2431
rect 7481 2397 7515 2431
rect 7941 2397 7975 2431
rect 9137 2397 9171 2431
rect 9229 2397 9263 2431
rect 9413 2397 9447 2431
rect 9597 2397 9631 2431
rect 10977 2397 11011 2431
rect 11529 2397 11563 2431
rect 11805 2397 11839 2431
rect 11897 2397 11931 2431
rect 12633 2397 12667 2431
rect 13461 2397 13495 2431
rect 14749 2397 14783 2431
rect 14841 2397 14875 2431
rect 2697 2329 2731 2363
rect 3893 2329 3927 2363
rect 4905 2329 4939 2363
rect 10241 2329 10275 2363
rect 14381 2329 14415 2363
rect 14473 2329 14507 2363
rect 6837 2261 6871 2295
rect 8953 2261 8987 2295
rect 10149 2261 10183 2295
<< metal1 >>
rect 1104 16346 15732 16368
rect 1104 16294 5858 16346
rect 5910 16294 5922 16346
rect 5974 16294 5986 16346
rect 6038 16294 6050 16346
rect 6102 16294 10734 16346
rect 10786 16294 10798 16346
rect 10850 16294 10862 16346
rect 10914 16294 10926 16346
rect 10978 16294 15732 16346
rect 1104 16272 15732 16294
rect 3878 16124 3884 16176
rect 3936 16164 3942 16176
rect 4893 16167 4951 16173
rect 4893 16164 4905 16167
rect 3936 16136 4905 16164
rect 3936 16124 3942 16136
rect 4893 16133 4905 16136
rect 4939 16133 4951 16167
rect 4893 16127 4951 16133
rect 7558 16124 7564 16176
rect 7616 16164 7622 16176
rect 7653 16167 7711 16173
rect 7653 16164 7665 16167
rect 7616 16136 7665 16164
rect 7616 16124 7622 16136
rect 7653 16133 7665 16136
rect 7699 16133 7711 16167
rect 7653 16127 7711 16133
rect 9674 16124 9680 16176
rect 9732 16164 9738 16176
rect 9953 16167 10011 16173
rect 9953 16164 9965 16167
rect 9732 16136 9965 16164
rect 9732 16124 9738 16136
rect 9953 16133 9965 16136
rect 9999 16133 10011 16167
rect 9953 16127 10011 16133
rect 13078 16124 13084 16176
rect 13136 16164 13142 16176
rect 13265 16167 13323 16173
rect 13265 16164 13277 16167
rect 13136 16136 13277 16164
rect 13136 16124 13142 16136
rect 13265 16133 13277 16136
rect 13311 16133 13323 16167
rect 16758 16164 16764 16176
rect 13265 16127 13323 16133
rect 14200 16136 16764 16164
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16056 1458 16108
rect 2866 16096 2872 16108
rect 2827 16068 2872 16096
rect 2866 16056 2872 16068
rect 2924 16056 2930 16108
rect 2958 16056 2964 16108
rect 3016 16096 3022 16108
rect 3234 16096 3240 16108
rect 3016 16068 3061 16096
rect 3195 16068 3240 16096
rect 3016 16056 3022 16068
rect 3234 16056 3240 16068
rect 3292 16056 3298 16108
rect 4246 16056 4252 16108
rect 4304 16096 4310 16108
rect 4341 16099 4399 16105
rect 4341 16096 4353 16099
rect 4304 16068 4353 16096
rect 4304 16056 4310 16068
rect 4341 16065 4353 16068
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16096 5135 16099
rect 5258 16096 5264 16108
rect 5123 16068 5264 16096
rect 5123 16065 5135 16068
rect 5077 16059 5135 16065
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 6365 16099 6423 16105
rect 6365 16096 6377 16099
rect 5776 16068 6377 16096
rect 5776 16056 5782 16068
rect 6365 16065 6377 16068
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 7837 16099 7895 16105
rect 7837 16065 7849 16099
rect 7883 16065 7895 16099
rect 9122 16096 9128 16108
rect 9083 16068 9128 16096
rect 7837 16059 7895 16065
rect 1673 16031 1731 16037
rect 1673 15997 1685 16031
rect 1719 16028 1731 16031
rect 6546 16028 6552 16040
rect 1719 16000 6552 16028
rect 1719 15997 1731 16000
rect 1673 15991 1731 15997
rect 6546 15988 6552 16000
rect 6604 15988 6610 16040
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 16028 6699 16031
rect 6822 16028 6828 16040
rect 6687 16000 6828 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 7852 16028 7880 16059
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 9214 16056 9220 16108
rect 9272 16096 9278 16108
rect 9493 16099 9551 16105
rect 9272 16068 9317 16096
rect 9272 16056 9278 16068
rect 9493 16065 9505 16099
rect 9539 16096 9551 16099
rect 9766 16096 9772 16108
rect 9539 16068 9772 16096
rect 9539 16065 9551 16068
rect 9493 16059 9551 16065
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 10134 16096 10140 16108
rect 10095 16068 10140 16096
rect 10134 16056 10140 16068
rect 10192 16056 10198 16108
rect 11238 16056 11244 16108
rect 11296 16096 11302 16108
rect 11517 16099 11575 16105
rect 11517 16096 11529 16099
rect 11296 16068 11529 16096
rect 11296 16056 11302 16068
rect 11517 16065 11529 16068
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16096 12587 16099
rect 14200 16096 14228 16136
rect 16758 16124 16764 16136
rect 16816 16124 16822 16176
rect 12575 16068 14228 16096
rect 14277 16099 14335 16105
rect 12575 16065 12587 16068
rect 12529 16059 12587 16065
rect 14277 16065 14289 16099
rect 14323 16096 14335 16099
rect 14550 16096 14556 16108
rect 14323 16068 14556 16096
rect 14323 16065 14335 16068
rect 14277 16059 14335 16065
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 14642 16056 14648 16108
rect 14700 16096 14706 16108
rect 14829 16099 14887 16105
rect 14829 16096 14841 16099
rect 14700 16068 14841 16096
rect 14700 16056 14706 16068
rect 14829 16065 14841 16068
rect 14875 16065 14887 16099
rect 15010 16096 15016 16108
rect 14971 16068 15016 16096
rect 14829 16059 14887 16065
rect 15010 16056 15016 16068
rect 15068 16056 15074 16108
rect 12618 16028 12624 16040
rect 7852 16000 12624 16028
rect 12618 15988 12624 16000
rect 12676 15988 12682 16040
rect 4154 15960 4160 15972
rect 4115 15932 4160 15960
rect 4154 15920 4160 15932
rect 4212 15920 4218 15972
rect 12713 15963 12771 15969
rect 12713 15929 12725 15963
rect 12759 15960 12771 15963
rect 13814 15960 13820 15972
rect 12759 15932 13820 15960
rect 12759 15929 12771 15932
rect 12713 15923 12771 15929
rect 13814 15920 13820 15932
rect 13872 15920 13878 15972
rect 2038 15852 2044 15904
rect 2096 15892 2102 15904
rect 2685 15895 2743 15901
rect 2685 15892 2697 15895
rect 2096 15864 2697 15892
rect 2096 15852 2102 15864
rect 2685 15861 2697 15864
rect 2731 15861 2743 15895
rect 3142 15892 3148 15904
rect 3103 15864 3148 15892
rect 2685 15855 2743 15861
rect 3142 15852 3148 15864
rect 3200 15852 3206 15904
rect 5442 15852 5448 15904
rect 5500 15892 5506 15904
rect 8941 15895 8999 15901
rect 8941 15892 8953 15895
rect 5500 15864 8953 15892
rect 5500 15852 5506 15864
rect 8941 15861 8953 15864
rect 8987 15861 8999 15895
rect 9398 15892 9404 15904
rect 9359 15864 9404 15892
rect 8941 15855 8999 15861
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 11698 15892 11704 15904
rect 11659 15864 11704 15892
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 12802 15852 12808 15904
rect 12860 15892 12866 15904
rect 13357 15895 13415 15901
rect 13357 15892 13369 15895
rect 12860 15864 13369 15892
rect 12860 15852 12866 15864
rect 13357 15861 13369 15864
rect 13403 15861 13415 15895
rect 13357 15855 13415 15861
rect 14093 15895 14151 15901
rect 14093 15861 14105 15895
rect 14139 15892 14151 15895
rect 14734 15892 14740 15904
rect 14139 15864 14740 15892
rect 14139 15861 14151 15864
rect 14093 15855 14151 15861
rect 14734 15852 14740 15864
rect 14792 15852 14798 15904
rect 1104 15802 15732 15824
rect 1104 15750 3420 15802
rect 3472 15750 3484 15802
rect 3536 15750 3548 15802
rect 3600 15750 3612 15802
rect 3664 15750 8296 15802
rect 8348 15750 8360 15802
rect 8412 15750 8424 15802
rect 8476 15750 8488 15802
rect 8540 15750 13172 15802
rect 13224 15750 13236 15802
rect 13288 15750 13300 15802
rect 13352 15750 13364 15802
rect 13416 15750 15732 15802
rect 1104 15728 15732 15750
rect 9214 15648 9220 15700
rect 9272 15688 9278 15700
rect 9401 15691 9459 15697
rect 9401 15688 9413 15691
rect 9272 15660 9413 15688
rect 9272 15648 9278 15660
rect 9401 15657 9413 15660
rect 9447 15657 9459 15691
rect 14642 15688 14648 15700
rect 14603 15660 14648 15688
rect 9401 15651 9459 15657
rect 14642 15648 14648 15660
rect 14700 15648 14706 15700
rect 2866 15580 2872 15632
rect 2924 15580 2930 15632
rect 5442 15620 5448 15632
rect 4816 15592 5448 15620
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15552 1547 15555
rect 1578 15552 1584 15564
rect 1535 15524 1584 15552
rect 1535 15521 1547 15524
rect 1489 15515 1547 15521
rect 1578 15512 1584 15524
rect 1636 15552 1642 15564
rect 2038 15552 2044 15564
rect 1636 15524 2044 15552
rect 1636 15512 1642 15524
rect 2038 15512 2044 15524
rect 2096 15512 2102 15564
rect 2685 15555 2743 15561
rect 2685 15521 2697 15555
rect 2731 15552 2743 15555
rect 2884 15552 2912 15580
rect 3237 15555 3295 15561
rect 3237 15552 3249 15555
rect 2731 15524 3249 15552
rect 2731 15521 2743 15524
rect 2685 15515 2743 15521
rect 3237 15521 3249 15524
rect 3283 15552 3295 15555
rect 4525 15555 4583 15561
rect 4525 15552 4537 15555
rect 3283 15524 4537 15552
rect 3283 15521 3295 15524
rect 3237 15515 3295 15521
rect 4525 15521 4537 15524
rect 4571 15521 4583 15555
rect 4816 15552 4844 15592
rect 5442 15580 5448 15592
rect 5500 15580 5506 15632
rect 8113 15623 8171 15629
rect 8113 15589 8125 15623
rect 8159 15589 8171 15623
rect 8113 15583 8171 15589
rect 11149 15623 11207 15629
rect 11149 15589 11161 15623
rect 11195 15589 11207 15623
rect 12894 15620 12900 15632
rect 12855 15592 12900 15620
rect 11149 15583 11207 15589
rect 4525 15515 4583 15521
rect 4724 15524 4844 15552
rect 4985 15555 5043 15561
rect 1670 15484 1676 15496
rect 1631 15456 1676 15484
rect 1670 15444 1676 15456
rect 1728 15484 1734 15496
rect 2869 15487 2927 15493
rect 1728 15456 1992 15484
rect 1728 15444 1734 15456
rect 1964 15425 1992 15456
rect 2869 15453 2881 15487
rect 2915 15484 2927 15487
rect 2958 15484 2964 15496
rect 2915 15456 2964 15484
rect 2915 15453 2927 15456
rect 2869 15447 2927 15453
rect 2958 15444 2964 15456
rect 3016 15484 3022 15496
rect 4724 15493 4752 15524
rect 4985 15521 4997 15555
rect 5031 15521 5043 15555
rect 4985 15515 5043 15521
rect 5721 15555 5779 15561
rect 5721 15521 5733 15555
rect 5767 15552 5779 15555
rect 8128 15552 8156 15583
rect 9398 15552 9404 15564
rect 5767 15524 6224 15552
rect 8128 15524 9404 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 4709 15487 4767 15493
rect 3016 15456 3188 15484
rect 3016 15444 3022 15456
rect 1949 15419 2007 15425
rect 1949 15385 1961 15419
rect 1995 15385 2007 15419
rect 1949 15379 2007 15385
rect 1854 15348 1860 15360
rect 1815 15320 1860 15348
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 2866 15308 2872 15360
rect 2924 15348 2930 15360
rect 3160 15357 3188 15456
rect 4709 15453 4721 15487
rect 4755 15453 4767 15487
rect 4709 15447 4767 15453
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15453 4859 15487
rect 4801 15447 4859 15453
rect 3053 15351 3111 15357
rect 3053 15348 3065 15351
rect 2924 15320 3065 15348
rect 2924 15308 2930 15320
rect 3053 15317 3065 15320
rect 3099 15317 3111 15351
rect 3053 15311 3111 15317
rect 3145 15351 3203 15357
rect 3145 15317 3157 15351
rect 3191 15348 3203 15351
rect 3418 15348 3424 15360
rect 3191 15320 3424 15348
rect 3191 15317 3203 15320
rect 3145 15311 3203 15317
rect 3418 15308 3424 15320
rect 3476 15308 3482 15360
rect 4816 15348 4844 15447
rect 5000 15416 5028 15515
rect 5077 15487 5135 15493
rect 5077 15453 5089 15487
rect 5123 15484 5135 15487
rect 5736 15484 5764 15515
rect 5123 15456 5764 15484
rect 5813 15487 5871 15493
rect 5123 15453 5135 15456
rect 5077 15447 5135 15453
rect 5813 15453 5825 15487
rect 5859 15453 5871 15487
rect 5813 15447 5871 15453
rect 5626 15416 5632 15428
rect 5000 15388 5632 15416
rect 5626 15376 5632 15388
rect 5684 15416 5690 15428
rect 5828 15416 5856 15447
rect 6196 15428 6224 15524
rect 9398 15512 9404 15524
rect 9456 15552 9462 15564
rect 9953 15555 10011 15561
rect 9953 15552 9965 15555
rect 9456 15524 9965 15552
rect 9456 15512 9462 15524
rect 7374 15444 7380 15496
rect 7432 15484 7438 15496
rect 7561 15487 7619 15493
rect 7561 15484 7573 15487
rect 7432 15456 7573 15484
rect 7432 15444 7438 15456
rect 7561 15453 7573 15456
rect 7607 15484 7619 15487
rect 7837 15487 7895 15493
rect 7837 15484 7849 15487
rect 7607 15456 7849 15484
rect 7607 15453 7619 15456
rect 7561 15447 7619 15453
rect 7837 15453 7849 15456
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 7926 15444 7932 15496
rect 7984 15484 7990 15496
rect 9692 15493 9720 15524
rect 9953 15521 9965 15524
rect 9999 15521 10011 15555
rect 11164 15552 11192 15583
rect 12894 15580 12900 15592
rect 12952 15580 12958 15632
rect 14921 15555 14979 15561
rect 14921 15552 14933 15555
rect 11164 15524 12020 15552
rect 9953 15515 10011 15521
rect 9585 15487 9643 15493
rect 7984 15456 8029 15484
rect 7984 15444 7990 15456
rect 9585 15453 9597 15487
rect 9631 15453 9643 15487
rect 9585 15447 9643 15453
rect 9677 15487 9735 15493
rect 9677 15453 9689 15487
rect 9723 15453 9735 15487
rect 9677 15447 9735 15453
rect 6089 15419 6147 15425
rect 6089 15416 6101 15419
rect 5684 15388 6101 15416
rect 5684 15376 5690 15388
rect 6089 15385 6101 15388
rect 6135 15385 6147 15419
rect 6089 15379 6147 15385
rect 6178 15376 6184 15428
rect 6236 15416 6242 15428
rect 7469 15419 7527 15425
rect 6236 15388 6281 15416
rect 6236 15376 6242 15388
rect 7469 15385 7481 15419
rect 7515 15416 7527 15419
rect 7944 15416 7972 15444
rect 7515 15388 7972 15416
rect 9600 15416 9628 15447
rect 10410 15444 10416 15496
rect 10468 15484 10474 15496
rect 10597 15487 10655 15493
rect 10597 15484 10609 15487
rect 10468 15456 10609 15484
rect 10468 15444 10474 15456
rect 10597 15453 10609 15456
rect 10643 15484 10655 15487
rect 10873 15487 10931 15493
rect 10873 15484 10885 15487
rect 10643 15456 10885 15484
rect 10643 15453 10655 15456
rect 10597 15447 10655 15453
rect 10873 15453 10885 15456
rect 10919 15453 10931 15487
rect 10873 15447 10931 15453
rect 10965 15487 11023 15493
rect 10965 15453 10977 15487
rect 11011 15453 11023 15487
rect 10965 15447 11023 15453
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15453 11667 15487
rect 11992 15484 12020 15524
rect 14384 15524 14933 15552
rect 12066 15484 12072 15496
rect 11979 15456 12072 15484
rect 11609 15447 11667 15453
rect 9766 15416 9772 15428
rect 9600 15388 9772 15416
rect 7515 15385 7527 15388
rect 7469 15379 7527 15385
rect 9766 15376 9772 15388
rect 9824 15416 9830 15428
rect 10045 15419 10103 15425
rect 10045 15416 10057 15419
rect 9824 15388 10057 15416
rect 9824 15376 9830 15388
rect 10045 15385 10057 15388
rect 10091 15416 10103 15419
rect 10318 15416 10324 15428
rect 10091 15388 10324 15416
rect 10091 15385 10103 15388
rect 10045 15379 10103 15385
rect 10318 15376 10324 15388
rect 10376 15376 10382 15428
rect 10502 15416 10508 15428
rect 10463 15388 10508 15416
rect 10502 15376 10508 15388
rect 10560 15416 10566 15428
rect 10980 15416 11008 15447
rect 10560 15388 11008 15416
rect 11624 15416 11652 15447
rect 12066 15444 12072 15456
rect 12124 15484 12130 15496
rect 12345 15487 12403 15493
rect 12345 15484 12357 15487
rect 12124 15456 12357 15484
rect 12124 15444 12130 15456
rect 12345 15453 12357 15456
rect 12391 15484 12403 15487
rect 12621 15487 12679 15493
rect 12621 15484 12633 15487
rect 12391 15456 12633 15484
rect 12391 15453 12403 15456
rect 12345 15447 12403 15453
rect 12621 15453 12633 15456
rect 12667 15453 12679 15487
rect 12621 15447 12679 15453
rect 12713 15487 12771 15493
rect 12713 15453 12725 15487
rect 12759 15453 12771 15487
rect 12713 15447 12771 15453
rect 12250 15416 12256 15428
rect 11624 15388 12020 15416
rect 12211 15388 12256 15416
rect 10560 15376 10566 15388
rect 5350 15348 5356 15360
rect 4816 15320 5356 15348
rect 5350 15308 5356 15320
rect 5408 15348 5414 15360
rect 5537 15351 5595 15357
rect 5537 15348 5549 15351
rect 5408 15320 5549 15348
rect 5408 15308 5414 15320
rect 5537 15317 5549 15320
rect 5583 15317 5595 15351
rect 11790 15348 11796 15360
rect 11751 15320 11796 15348
rect 5537 15311 5595 15317
rect 11790 15308 11796 15320
rect 11848 15308 11854 15360
rect 11992 15348 12020 15388
rect 12250 15376 12256 15388
rect 12308 15416 12314 15428
rect 12728 15416 12756 15447
rect 12986 15444 12992 15496
rect 13044 15484 13050 15496
rect 13357 15487 13415 15493
rect 13357 15484 13369 15487
rect 13044 15456 13369 15484
rect 13044 15444 13050 15456
rect 13357 15453 13369 15456
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15484 13599 15487
rect 14182 15484 14188 15496
rect 13587 15456 14188 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 14182 15444 14188 15456
rect 14240 15444 14246 15496
rect 14274 15444 14280 15496
rect 14332 15484 14338 15496
rect 14384 15493 14412 15524
rect 14921 15521 14933 15524
rect 14967 15521 14979 15555
rect 14921 15515 14979 15521
rect 14369 15487 14427 15493
rect 14369 15484 14381 15487
rect 14332 15456 14381 15484
rect 14332 15444 14338 15456
rect 14369 15453 14381 15456
rect 14415 15453 14427 15487
rect 14737 15487 14795 15493
rect 14737 15484 14749 15487
rect 14369 15447 14427 15453
rect 14476 15456 14749 15484
rect 14476 15428 14504 15456
rect 14737 15453 14749 15456
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 14458 15416 14464 15428
rect 12308 15388 12756 15416
rect 12820 15388 14320 15416
rect 14371 15388 14464 15416
rect 12308 15376 12314 15388
rect 12820 15348 12848 15388
rect 11992 15320 12848 15348
rect 13449 15351 13507 15357
rect 13449 15317 13461 15351
rect 13495 15348 13507 15351
rect 13998 15348 14004 15360
rect 13495 15320 14004 15348
rect 13495 15317 13507 15320
rect 13449 15311 13507 15317
rect 13998 15308 14004 15320
rect 14056 15308 14062 15360
rect 14292 15348 14320 15388
rect 14458 15376 14464 15388
rect 14516 15376 14522 15428
rect 14918 15348 14924 15360
rect 14292 15320 14924 15348
rect 14918 15308 14924 15320
rect 14976 15308 14982 15360
rect 1104 15258 15732 15280
rect 1104 15206 5858 15258
rect 5910 15206 5922 15258
rect 5974 15206 5986 15258
rect 6038 15206 6050 15258
rect 6102 15206 10734 15258
rect 10786 15206 10798 15258
rect 10850 15206 10862 15258
rect 10914 15206 10926 15258
rect 10978 15206 15732 15258
rect 1104 15184 15732 15206
rect 1946 15104 1952 15156
rect 2004 15144 2010 15156
rect 2501 15147 2559 15153
rect 2501 15144 2513 15147
rect 2004 15116 2513 15144
rect 2004 15104 2010 15116
rect 2501 15113 2513 15116
rect 2547 15113 2559 15147
rect 3418 15144 3424 15156
rect 3379 15116 3424 15144
rect 2501 15107 2559 15113
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 5350 15144 5356 15156
rect 5311 15116 5356 15144
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 6178 15104 6184 15156
rect 6236 15144 6242 15156
rect 7101 15147 7159 15153
rect 7101 15144 7113 15147
rect 6236 15116 7113 15144
rect 6236 15104 6242 15116
rect 7101 15113 7113 15116
rect 7147 15113 7159 15147
rect 7101 15107 7159 15113
rect 9214 15104 9220 15156
rect 9272 15144 9278 15156
rect 9309 15147 9367 15153
rect 9309 15144 9321 15147
rect 9272 15116 9321 15144
rect 9272 15104 9278 15116
rect 9309 15113 9321 15116
rect 9355 15113 9367 15147
rect 9309 15107 9367 15113
rect 9401 15147 9459 15153
rect 9401 15113 9413 15147
rect 9447 15144 9459 15147
rect 10134 15144 10140 15156
rect 9447 15116 10140 15144
rect 9447 15113 9459 15116
rect 9401 15107 9459 15113
rect 1854 15036 1860 15088
rect 1912 15076 1918 15088
rect 2593 15079 2651 15085
rect 2593 15076 2605 15079
rect 1912 15048 2605 15076
rect 1912 15036 1918 15048
rect 2593 15045 2605 15048
rect 2639 15045 2651 15079
rect 2593 15039 2651 15045
rect 1578 15008 1584 15020
rect 1539 14980 1584 15008
rect 1578 14968 1584 14980
rect 1636 14968 1642 15020
rect 1670 14968 1676 15020
rect 1728 15008 1734 15020
rect 1949 15011 2007 15017
rect 1728 14980 1773 15008
rect 1728 14968 1734 14980
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 2038 15008 2044 15020
rect 1995 14980 2044 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2038 14968 2044 14980
rect 2096 14968 2102 15020
rect 3142 14968 3148 15020
rect 3200 15008 3206 15020
rect 3697 15011 3755 15017
rect 3697 15008 3709 15011
rect 3200 14980 3709 15008
rect 3200 14968 3206 14980
rect 3697 14977 3709 14980
rect 3743 15008 3755 15011
rect 3973 15011 4031 15017
rect 3973 15008 3985 15011
rect 3743 14980 3985 15008
rect 3743 14977 3755 14980
rect 3697 14971 3755 14977
rect 3973 14977 3985 14980
rect 4019 14977 4031 15011
rect 5368 15008 5396 15104
rect 7926 15076 7932 15088
rect 7300 15048 7932 15076
rect 7300 15017 7328 15048
rect 7926 15036 7932 15048
rect 7984 15036 7990 15088
rect 5629 15011 5687 15017
rect 5629 15008 5641 15011
rect 5368 14980 5641 15008
rect 3973 14971 4031 14977
rect 5629 14977 5641 14980
rect 5675 14977 5687 15011
rect 5629 14971 5687 14977
rect 7285 15011 7343 15017
rect 7285 14977 7297 15011
rect 7331 14977 7343 15011
rect 7285 14971 7343 14977
rect 7374 14968 7380 15020
rect 7432 15008 7438 15020
rect 7650 15008 7656 15020
rect 7432 14980 7477 15008
rect 7611 14980 7656 15008
rect 7432 14968 7438 14980
rect 7650 14968 7656 14980
rect 7708 14968 7714 15020
rect 9324 15008 9352 15107
rect 10134 15104 10140 15116
rect 10192 15104 10198 15156
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12897 15147 12955 15153
rect 12897 15144 12909 15147
rect 12676 15116 12909 15144
rect 12676 15104 12682 15116
rect 12897 15113 12909 15116
rect 12943 15113 12955 15147
rect 14458 15144 14464 15156
rect 14419 15116 14464 15144
rect 12897 15107 12955 15113
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 12805 15079 12863 15085
rect 12805 15076 12817 15079
rect 11900 15048 12817 15076
rect 11900 15017 11928 15048
rect 12805 15045 12817 15048
rect 12851 15045 12863 15079
rect 12805 15039 12863 15045
rect 9585 15011 9643 15017
rect 9585 15008 9597 15011
rect 9324 14980 9597 15008
rect 9585 14977 9597 14980
rect 9631 14977 9643 15011
rect 9585 14971 9643 14977
rect 9769 15011 9827 15017
rect 9769 14977 9781 15011
rect 9815 15008 9827 15011
rect 11609 15011 11667 15017
rect 11609 15008 11621 15011
rect 9815 14980 11621 15008
rect 9815 14977 9827 14980
rect 9769 14971 9827 14977
rect 11609 14977 11621 14980
rect 11655 14977 11667 15011
rect 11609 14971 11667 14977
rect 11793 15011 11851 15017
rect 11793 14977 11805 15011
rect 11839 14977 11851 15011
rect 11793 14971 11851 14977
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 14977 11943 15011
rect 11885 14971 11943 14977
rect 12161 15011 12219 15017
rect 12161 14977 12173 15011
rect 12207 15008 12219 15011
rect 12250 15008 12256 15020
rect 12207 14980 12256 15008
rect 12207 14977 12219 14980
rect 12161 14971 12219 14977
rect 3234 14900 3240 14952
rect 3292 14940 3298 14952
rect 3605 14943 3663 14949
rect 3605 14940 3617 14943
rect 3292 14912 3617 14940
rect 3292 14900 3298 14912
rect 3605 14909 3617 14912
rect 3651 14940 3663 14943
rect 4062 14940 4068 14952
rect 3651 14912 4068 14940
rect 3651 14909 3663 14912
rect 3605 14903 3663 14909
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 5261 14943 5319 14949
rect 5261 14909 5273 14943
rect 5307 14940 5319 14943
rect 5442 14940 5448 14952
rect 5307 14912 5448 14940
rect 5307 14909 5319 14912
rect 5261 14903 5319 14909
rect 5442 14900 5448 14912
rect 5500 14940 5506 14952
rect 5813 14943 5871 14949
rect 5813 14940 5825 14943
rect 5500 14912 5825 14940
rect 5500 14900 5506 14912
rect 5813 14909 5825 14912
rect 5859 14909 5871 14943
rect 5813 14903 5871 14909
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 9217 14943 9275 14949
rect 9217 14940 9229 14943
rect 9180 14912 9229 14940
rect 9180 14900 9186 14912
rect 9217 14909 9229 14912
rect 9263 14940 9275 14943
rect 9784 14940 9812 14971
rect 9263 14912 9812 14940
rect 9263 14909 9275 14912
rect 9217 14903 9275 14909
rect 14 14832 20 14884
rect 72 14872 78 14884
rect 4154 14872 4160 14884
rect 72 14844 4160 14872
rect 72 14832 78 14844
rect 4154 14832 4160 14844
rect 4212 14832 4218 14884
rect 11808 14872 11836 14971
rect 12250 14968 12256 14980
rect 12308 14968 12314 15020
rect 12820 15008 12848 15039
rect 12894 15008 12900 15020
rect 12807 14980 12900 15008
rect 12894 14968 12900 14980
rect 12952 15008 12958 15020
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 12952 14980 13093 15008
rect 12952 14968 12958 14980
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 12066 14940 12072 14952
rect 12027 14912 12072 14940
rect 12066 14900 12072 14912
rect 12124 14900 12130 14952
rect 12713 14943 12771 14949
rect 12713 14909 12725 14943
rect 12759 14940 12771 14943
rect 13265 14943 13323 14949
rect 13265 14940 13277 14943
rect 12759 14912 13277 14940
rect 12759 14909 12771 14912
rect 12713 14903 12771 14909
rect 13265 14909 13277 14912
rect 13311 14940 13323 14943
rect 13538 14940 13544 14952
rect 13311 14912 13544 14940
rect 13311 14909 13323 14912
rect 13265 14903 13323 14909
rect 12728 14872 12756 14903
rect 13538 14900 13544 14912
rect 13596 14900 13602 14952
rect 13722 14900 13728 14952
rect 13780 14940 13786 14952
rect 13817 14943 13875 14949
rect 13817 14940 13829 14943
rect 13780 14912 13829 14940
rect 13780 14900 13786 14912
rect 13817 14909 13829 14912
rect 13863 14909 13875 14943
rect 13817 14903 13875 14909
rect 11808 14844 12756 14872
rect 13832 14872 13860 14903
rect 13906 14900 13912 14952
rect 13964 14940 13970 14952
rect 14200 14940 14228 14971
rect 13964 14912 14228 14940
rect 14277 14943 14335 14949
rect 13964 14900 13970 14912
rect 14277 14909 14289 14943
rect 14323 14909 14335 14943
rect 14277 14903 14335 14909
rect 14292 14872 14320 14903
rect 13832 14844 14320 14872
rect 1397 14807 1455 14813
rect 1397 14773 1409 14807
rect 1443 14804 1455 14807
rect 1578 14804 1584 14816
rect 1443 14776 1584 14804
rect 1443 14773 1455 14776
rect 1397 14767 1455 14773
rect 1578 14764 1584 14776
rect 1636 14764 1642 14816
rect 1857 14807 1915 14813
rect 1857 14773 1869 14807
rect 1903 14804 1915 14807
rect 2222 14804 2228 14816
rect 1903 14776 2228 14804
rect 1903 14773 1915 14776
rect 1857 14767 1915 14773
rect 2222 14764 2228 14776
rect 2280 14764 2286 14816
rect 5537 14807 5595 14813
rect 5537 14773 5549 14807
rect 5583 14804 5595 14807
rect 6638 14804 6644 14816
rect 5583 14776 6644 14804
rect 5583 14773 5595 14776
rect 5537 14767 5595 14773
rect 6638 14764 6644 14776
rect 6696 14764 6702 14816
rect 7558 14804 7564 14816
rect 7519 14776 7564 14804
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 1104 14714 15732 14736
rect 1104 14662 3420 14714
rect 3472 14662 3484 14714
rect 3536 14662 3548 14714
rect 3600 14662 3612 14714
rect 3664 14662 8296 14714
rect 8348 14662 8360 14714
rect 8412 14662 8424 14714
rect 8476 14662 8488 14714
rect 8540 14662 13172 14714
rect 13224 14662 13236 14714
rect 13288 14662 13300 14714
rect 13352 14662 13364 14714
rect 13416 14662 15732 14714
rect 1104 14640 15732 14662
rect 1670 14600 1676 14612
rect 1631 14572 1676 14600
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 4525 14603 4583 14609
rect 4525 14600 4537 14603
rect 4120 14572 4537 14600
rect 4120 14560 4126 14572
rect 4525 14569 4537 14572
rect 4571 14569 4583 14603
rect 4525 14563 4583 14569
rect 7009 14603 7067 14609
rect 7009 14569 7021 14603
rect 7055 14600 7067 14603
rect 7374 14600 7380 14612
rect 7055 14572 7380 14600
rect 7055 14569 7067 14572
rect 7009 14563 7067 14569
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 7926 14560 7932 14612
rect 7984 14600 7990 14612
rect 8941 14603 8999 14609
rect 8941 14600 8953 14603
rect 7984 14572 8953 14600
rect 7984 14560 7990 14572
rect 8941 14569 8953 14572
rect 8987 14569 8999 14603
rect 10410 14600 10416 14612
rect 10371 14572 10416 14600
rect 8941 14563 8999 14569
rect 10410 14560 10416 14572
rect 10468 14560 10474 14612
rect 12250 14560 12256 14612
rect 12308 14600 12314 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 12308 14572 13001 14600
rect 12308 14560 12314 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13596 14572 14105 14600
rect 13596 14560 13602 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 14093 14563 14151 14569
rect 4985 14535 5043 14541
rect 4985 14501 4997 14535
rect 5031 14532 5043 14535
rect 5074 14532 5080 14544
rect 5031 14504 5080 14532
rect 5031 14501 5043 14504
rect 4985 14495 5043 14501
rect 5074 14492 5080 14504
rect 5132 14492 5138 14544
rect 7650 14532 7656 14544
rect 7208 14504 7656 14532
rect 1857 14467 1915 14473
rect 1857 14433 1869 14467
rect 1903 14464 1915 14467
rect 2038 14464 2044 14476
rect 1903 14436 2044 14464
rect 1903 14433 1915 14436
rect 1857 14427 1915 14433
rect 2038 14424 2044 14436
rect 2096 14464 2102 14476
rect 7208 14473 7236 14504
rect 7650 14492 7656 14504
rect 7708 14532 7714 14544
rect 7708 14504 7788 14532
rect 7708 14492 7714 14504
rect 7193 14467 7251 14473
rect 2096 14436 2360 14464
rect 2096 14424 2102 14436
rect 1949 14399 2007 14405
rect 1949 14365 1961 14399
rect 1995 14396 2007 14399
rect 1995 14368 2268 14396
rect 1995 14365 2007 14368
rect 1949 14359 2007 14365
rect 2240 14340 2268 14368
rect 2222 14328 2228 14340
rect 2183 14300 2228 14328
rect 2222 14288 2228 14300
rect 2280 14288 2286 14340
rect 2332 14337 2360 14436
rect 7193 14433 7205 14467
rect 7239 14433 7251 14467
rect 7193 14427 7251 14433
rect 4706 14396 4712 14408
rect 4667 14368 4712 14396
rect 4706 14356 4712 14368
rect 4764 14356 4770 14408
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 5077 14399 5135 14405
rect 4856 14368 4901 14396
rect 4856 14356 4862 14368
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5534 14396 5540 14408
rect 5123 14368 5540 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 7285 14399 7343 14405
rect 7285 14365 7297 14399
rect 7331 14396 7343 14399
rect 7653 14399 7711 14405
rect 7331 14368 7604 14396
rect 7331 14365 7343 14368
rect 7285 14359 7343 14365
rect 7576 14340 7604 14368
rect 7653 14365 7665 14399
rect 7699 14395 7711 14399
rect 7760 14396 7788 14504
rect 9646 14504 11192 14532
rect 9646 14464 9674 14504
rect 8036 14436 9674 14464
rect 10597 14467 10655 14473
rect 8036 14396 8064 14436
rect 10597 14433 10609 14467
rect 10643 14464 10655 14467
rect 11164 14464 11192 14504
rect 12434 14492 12440 14544
rect 12492 14532 12498 14544
rect 12529 14535 12587 14541
rect 12529 14532 12541 14535
rect 12492 14504 12541 14532
rect 12492 14492 12498 14504
rect 12529 14501 12541 14504
rect 12575 14501 12587 14535
rect 12529 14495 12587 14501
rect 13906 14492 13912 14544
rect 13964 14532 13970 14544
rect 14553 14535 14611 14541
rect 14553 14532 14565 14535
rect 13964 14504 14565 14532
rect 13964 14492 13970 14504
rect 14553 14501 14565 14504
rect 14599 14501 14611 14535
rect 14553 14495 14611 14501
rect 12618 14464 12624 14476
rect 10643 14436 11100 14464
rect 11164 14436 12624 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 7760 14395 8064 14396
rect 7699 14368 8064 14395
rect 8297 14399 8355 14405
rect 7699 14367 7788 14368
rect 7699 14365 7711 14367
rect 7653 14359 7711 14365
rect 8297 14365 8309 14399
rect 8343 14365 8355 14399
rect 8297 14359 8355 14365
rect 2317 14331 2375 14337
rect 2317 14297 2329 14331
rect 2363 14328 2375 14331
rect 2682 14328 2688 14340
rect 2363 14300 2688 14328
rect 2363 14297 2375 14300
rect 2317 14291 2375 14297
rect 2682 14288 2688 14300
rect 2740 14288 2746 14340
rect 7558 14328 7564 14340
rect 7519 14300 7564 14328
rect 7558 14288 7564 14300
rect 7616 14288 7622 14340
rect 8312 14328 8340 14359
rect 9858 14356 9864 14408
rect 9916 14396 9922 14408
rect 9953 14399 10011 14405
rect 9953 14396 9965 14399
rect 9916 14368 9965 14396
rect 9916 14356 9922 14368
rect 9953 14365 9965 14368
rect 9999 14365 10011 14399
rect 9953 14359 10011 14365
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14396 10747 14399
rect 10735 14368 11008 14396
rect 10735 14365 10747 14368
rect 10689 14359 10747 14365
rect 7668 14300 8340 14328
rect 9125 14331 9183 14337
rect 4890 14220 4896 14272
rect 4948 14260 4954 14272
rect 7282 14260 7288 14272
rect 4948 14232 7288 14260
rect 4948 14220 4954 14232
rect 7282 14220 7288 14232
rect 7340 14260 7346 14272
rect 7668 14260 7696 14300
rect 9125 14297 9137 14331
rect 9171 14297 9183 14331
rect 9125 14291 9183 14297
rect 9309 14331 9367 14337
rect 9309 14297 9321 14331
rect 9355 14328 9367 14331
rect 9582 14328 9588 14340
rect 9355 14300 9588 14328
rect 9355 14297 9367 14300
rect 9309 14291 9367 14297
rect 7340 14232 7696 14260
rect 7340 14220 7346 14232
rect 8110 14220 8116 14272
rect 8168 14260 8174 14272
rect 8205 14263 8263 14269
rect 8205 14260 8217 14263
rect 8168 14232 8217 14260
rect 8168 14220 8174 14232
rect 8205 14229 8217 14232
rect 8251 14229 8263 14263
rect 9140 14260 9168 14291
rect 9582 14288 9588 14300
rect 9640 14288 9646 14340
rect 10980 14337 11008 14368
rect 11072 14340 11100 14436
rect 12618 14424 12624 14436
rect 12676 14424 12682 14476
rect 13722 14424 13728 14476
rect 13780 14464 13786 14476
rect 13780 14436 14688 14464
rect 13780 14424 13786 14436
rect 11790 14396 11796 14408
rect 11703 14368 11796 14396
rect 11790 14356 11796 14368
rect 11848 14396 11854 14408
rect 12066 14396 12072 14408
rect 11848 14368 12072 14396
rect 11848 14356 11854 14368
rect 12066 14356 12072 14368
rect 12124 14356 12130 14408
rect 12158 14356 12164 14408
rect 12216 14396 12222 14408
rect 12437 14399 12495 14405
rect 12437 14396 12449 14399
rect 12216 14368 12449 14396
rect 12216 14356 12222 14368
rect 12437 14365 12449 14368
rect 12483 14365 12495 14399
rect 12710 14396 12716 14408
rect 12671 14368 12716 14396
rect 12437 14359 12495 14365
rect 12710 14356 12716 14368
rect 12768 14356 12774 14408
rect 12802 14356 12808 14408
rect 12860 14396 12866 14408
rect 14274 14396 14280 14408
rect 12860 14368 12905 14396
rect 14187 14368 14280 14396
rect 12860 14356 12866 14368
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14396 14427 14399
rect 14458 14396 14464 14408
rect 14415 14368 14464 14396
rect 14415 14365 14427 14368
rect 14369 14359 14427 14365
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 14660 14405 14688 14436
rect 14645 14399 14703 14405
rect 14645 14365 14657 14399
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 10965 14331 11023 14337
rect 10965 14297 10977 14331
rect 11011 14297 11023 14331
rect 10965 14291 11023 14297
rect 9398 14260 9404 14272
rect 9140 14232 9404 14260
rect 8205 14223 8263 14229
rect 9398 14220 9404 14232
rect 9456 14260 9462 14272
rect 9769 14263 9827 14269
rect 9769 14260 9781 14263
rect 9456 14232 9781 14260
rect 9456 14220 9462 14232
rect 9769 14229 9781 14232
rect 9815 14229 9827 14263
rect 10980 14260 11008 14291
rect 11054 14288 11060 14340
rect 11112 14328 11118 14340
rect 14292 14328 14320 14356
rect 14734 14328 14740 14340
rect 11112 14300 11157 14328
rect 14292 14300 14740 14328
rect 11112 14288 11118 14300
rect 14734 14288 14740 14300
rect 14792 14288 14798 14340
rect 11146 14260 11152 14272
rect 10980 14232 11152 14260
rect 9769 14223 9827 14229
rect 11146 14220 11152 14232
rect 11204 14220 11210 14272
rect 11885 14263 11943 14269
rect 11885 14229 11897 14263
rect 11931 14260 11943 14263
rect 14366 14260 14372 14272
rect 11931 14232 14372 14260
rect 11931 14229 11943 14232
rect 11885 14223 11943 14229
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 1104 14170 15732 14192
rect 1104 14118 5858 14170
rect 5910 14118 5922 14170
rect 5974 14118 5986 14170
rect 6038 14118 6050 14170
rect 6102 14118 10734 14170
rect 10786 14118 10798 14170
rect 10850 14118 10862 14170
rect 10914 14118 10926 14170
rect 10978 14118 15732 14170
rect 1104 14096 15732 14118
rect 3142 14056 3148 14068
rect 3103 14028 3148 14056
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 4798 14056 4804 14068
rect 4759 14028 4804 14056
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 7558 14016 7564 14068
rect 7616 14056 7622 14068
rect 7837 14059 7895 14065
rect 7837 14056 7849 14059
rect 7616 14028 7849 14056
rect 7616 14016 7622 14028
rect 7837 14025 7849 14028
rect 7883 14025 7895 14059
rect 10318 14056 10324 14068
rect 10279 14028 10324 14056
rect 7837 14019 7895 14025
rect 10318 14016 10324 14028
rect 10376 14016 10382 14068
rect 13449 14059 13507 14065
rect 12406 14028 13308 14056
rect 2041 13991 2099 13997
rect 2041 13957 2053 13991
rect 2087 13988 2099 13991
rect 4890 13988 4896 14000
rect 2087 13960 4896 13988
rect 2087 13957 2099 13960
rect 2041 13951 2099 13957
rect 4890 13948 4896 13960
rect 4948 13948 4954 14000
rect 9306 13948 9312 14000
rect 9364 13988 9370 14000
rect 9677 13991 9735 13997
rect 9677 13988 9689 13991
rect 9364 13960 9689 13988
rect 9364 13948 9370 13960
rect 9677 13957 9689 13960
rect 9723 13957 9735 13991
rect 9677 13951 9735 13957
rect 10410 13948 10416 14000
rect 10468 13988 10474 14000
rect 11146 13988 11152 14000
rect 10468 13960 10640 13988
rect 11059 13960 11152 13988
rect 10468 13948 10474 13960
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 2406 13880 2412 13932
rect 2464 13920 2470 13932
rect 2593 13923 2651 13929
rect 2593 13920 2605 13923
rect 2464 13892 2605 13920
rect 2464 13880 2470 13892
rect 2593 13889 2605 13892
rect 2639 13920 2651 13923
rect 2869 13923 2927 13929
rect 2869 13920 2881 13923
rect 2639 13892 2881 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 2869 13889 2881 13892
rect 2915 13889 2927 13923
rect 5074 13920 5080 13932
rect 5035 13892 5080 13920
rect 2869 13883 2927 13889
rect 5074 13880 5080 13892
rect 5132 13920 5138 13932
rect 5353 13923 5411 13929
rect 5353 13920 5365 13923
rect 5132 13892 5365 13920
rect 5132 13880 5138 13892
rect 5353 13889 5365 13892
rect 5399 13889 5411 13923
rect 5353 13883 5411 13889
rect 5718 13880 5724 13932
rect 5776 13920 5782 13932
rect 6730 13920 6736 13932
rect 5776 13892 6736 13920
rect 5776 13880 5782 13892
rect 6730 13880 6736 13892
rect 6788 13920 6794 13932
rect 6917 13923 6975 13929
rect 6917 13920 6929 13923
rect 6788 13892 6929 13920
rect 6788 13880 6794 13892
rect 6917 13889 6929 13892
rect 6963 13889 6975 13923
rect 6917 13883 6975 13889
rect 8113 13923 8171 13929
rect 8113 13889 8125 13923
rect 8159 13920 8171 13923
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 8159 13892 8401 13920
rect 8159 13889 8171 13892
rect 8113 13883 8171 13889
rect 8389 13889 8401 13892
rect 8435 13920 8447 13923
rect 8938 13920 8944 13932
rect 8435 13892 8944 13920
rect 8435 13889 8447 13892
rect 8389 13883 8447 13889
rect 8938 13880 8944 13892
rect 8996 13880 9002 13932
rect 9490 13920 9496 13932
rect 9451 13892 9496 13920
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 9861 13923 9919 13929
rect 9861 13889 9873 13923
rect 9907 13920 9919 13923
rect 10502 13920 10508 13932
rect 9907 13892 10508 13920
rect 9907 13889 9919 13892
rect 9861 13883 9919 13889
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 10612 13929 10640 13960
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13889 10655 13923
rect 10870 13920 10876 13932
rect 10831 13892 10876 13920
rect 10597 13883 10655 13889
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13852 2559 13855
rect 2961 13855 3019 13861
rect 2961 13852 2973 13855
rect 2547 13824 2973 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 2961 13821 2973 13824
rect 3007 13852 3019 13855
rect 3142 13852 3148 13864
rect 3007 13824 3148 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 3142 13812 3148 13824
rect 3200 13812 3206 13864
rect 4985 13855 5043 13861
rect 4985 13821 4997 13855
rect 5031 13852 5043 13855
rect 5445 13855 5503 13861
rect 5445 13852 5457 13855
rect 5031 13824 5457 13852
rect 5031 13821 5043 13824
rect 4985 13815 5043 13821
rect 5445 13821 5457 13824
rect 5491 13852 5503 13855
rect 5534 13852 5540 13864
rect 5491 13824 5540 13852
rect 5491 13821 5503 13824
rect 5445 13815 5503 13821
rect 5534 13812 5540 13824
rect 5592 13852 5598 13864
rect 5810 13852 5816 13864
rect 5592 13824 5816 13852
rect 5592 13812 5598 13824
rect 5810 13812 5816 13824
rect 5868 13812 5874 13864
rect 8018 13852 8024 13864
rect 7979 13824 8024 13852
rect 8018 13812 8024 13824
rect 8076 13852 8082 13864
rect 8481 13855 8539 13861
rect 8481 13852 8493 13855
rect 8076 13824 8493 13852
rect 8076 13812 8082 13824
rect 8481 13821 8493 13824
rect 8527 13821 8539 13855
rect 8481 13815 8539 13821
rect 10781 13855 10839 13861
rect 10781 13821 10793 13855
rect 10827 13852 10839 13855
rect 11072 13852 11100 13960
rect 11146 13948 11152 13960
rect 11204 13988 11210 14000
rect 12406 13988 12434 14028
rect 12710 13988 12716 14000
rect 11204 13960 12434 13988
rect 12623 13960 12716 13988
rect 11204 13948 11210 13960
rect 11698 13920 11704 13932
rect 11659 13892 11704 13920
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13920 12219 13923
rect 12250 13920 12256 13932
rect 12207 13892 12256 13920
rect 12207 13889 12219 13892
rect 12161 13883 12219 13889
rect 12250 13880 12256 13892
rect 12308 13880 12314 13932
rect 10827 13824 11100 13852
rect 10827 13821 10839 13824
rect 10781 13815 10839 13821
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 12636 13852 12664 13960
rect 12710 13948 12716 13960
rect 12768 13988 12774 14000
rect 13280 13988 13308 14028
rect 13449 14025 13461 14059
rect 13495 14056 13507 14059
rect 13906 14056 13912 14068
rect 13495 14028 13912 14056
rect 13495 14025 13507 14028
rect 13449 14019 13507 14025
rect 13906 14016 13912 14028
rect 13964 14016 13970 14068
rect 12768 13960 13216 13988
rect 13280 13960 13676 13988
rect 12768 13948 12774 13960
rect 12802 13920 12808 13932
rect 12715 13892 12808 13920
rect 12802 13880 12808 13892
rect 12860 13920 12866 13932
rect 13188 13929 13216 13960
rect 13173 13923 13231 13929
rect 12860 13892 13124 13920
rect 12860 13880 12866 13892
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12584 13824 12909 13852
rect 12584 13812 12590 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 13096 13852 13124 13892
rect 13173 13889 13185 13923
rect 13219 13889 13231 13923
rect 13173 13883 13231 13889
rect 13265 13855 13323 13861
rect 13265 13852 13277 13855
rect 13096 13824 13277 13852
rect 12897 13815 12955 13821
rect 13265 13821 13277 13824
rect 13311 13852 13323 13855
rect 13538 13852 13544 13864
rect 13311 13824 13544 13852
rect 13311 13821 13323 13824
rect 13265 13815 13323 13821
rect 13538 13812 13544 13824
rect 13596 13812 13602 13864
rect 13648 13852 13676 13960
rect 13814 13880 13820 13932
rect 13872 13920 13878 13932
rect 14093 13923 14151 13929
rect 14093 13920 14105 13923
rect 13872 13892 14105 13920
rect 13872 13880 13878 13892
rect 14093 13889 14105 13892
rect 14139 13889 14151 13923
rect 14826 13920 14832 13932
rect 14787 13892 14832 13920
rect 14093 13883 14151 13889
rect 14826 13880 14832 13892
rect 14884 13880 14890 13932
rect 13906 13852 13912 13864
rect 13648 13824 13912 13852
rect 13906 13812 13912 13824
rect 13964 13812 13970 13864
rect 14185 13855 14243 13861
rect 14185 13852 14197 13855
rect 14016 13824 14197 13852
rect 6178 13744 6184 13796
rect 6236 13784 6242 13796
rect 12802 13784 12808 13796
rect 6236 13756 12808 13784
rect 6236 13744 6242 13756
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 13630 13744 13636 13796
rect 13688 13784 13694 13796
rect 14016 13784 14044 13824
rect 14185 13821 14197 13824
rect 14231 13821 14243 13855
rect 15010 13852 15016 13864
rect 14971 13824 15016 13852
rect 14185 13815 14243 13821
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 13688 13756 14044 13784
rect 13688 13744 13694 13756
rect 7098 13716 7104 13728
rect 7059 13688 7104 13716
rect 7098 13676 7104 13688
rect 7156 13676 7162 13728
rect 11054 13676 11060 13728
rect 11112 13716 11118 13728
rect 11609 13719 11667 13725
rect 11609 13716 11621 13719
rect 11112 13688 11621 13716
rect 11112 13676 11118 13688
rect 11609 13685 11621 13688
rect 11655 13685 11667 13719
rect 11609 13679 11667 13685
rect 12345 13719 12403 13725
rect 12345 13685 12357 13719
rect 12391 13716 12403 13719
rect 12618 13716 12624 13728
rect 12391 13688 12624 13716
rect 12391 13685 12403 13688
rect 12345 13679 12403 13685
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 12820 13716 12848 13744
rect 15102 13716 15108 13728
rect 12820 13688 15108 13716
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 1104 13626 15732 13648
rect 1104 13574 3420 13626
rect 3472 13574 3484 13626
rect 3536 13574 3548 13626
rect 3600 13574 3612 13626
rect 3664 13574 8296 13626
rect 8348 13574 8360 13626
rect 8412 13574 8424 13626
rect 8476 13574 8488 13626
rect 8540 13574 13172 13626
rect 13224 13574 13236 13626
rect 13288 13574 13300 13626
rect 13352 13574 13364 13626
rect 13416 13574 15732 13626
rect 1104 13552 15732 13574
rect 2682 13512 2688 13524
rect 2643 13484 2688 13512
rect 2682 13472 2688 13484
rect 2740 13472 2746 13524
rect 5537 13515 5595 13521
rect 5537 13481 5549 13515
rect 5583 13512 5595 13515
rect 5626 13512 5632 13524
rect 5583 13484 5632 13512
rect 5583 13481 5595 13484
rect 5537 13475 5595 13481
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 7190 13512 7196 13524
rect 7151 13484 7196 13512
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7377 13515 7435 13521
rect 7377 13481 7389 13515
rect 7423 13512 7435 13515
rect 8018 13512 8024 13524
rect 7423 13484 8024 13512
rect 7423 13481 7435 13484
rect 7377 13475 7435 13481
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 8938 13512 8944 13524
rect 8899 13484 8944 13512
rect 8938 13472 8944 13484
rect 8996 13472 9002 13524
rect 11149 13515 11207 13521
rect 11149 13481 11161 13515
rect 11195 13512 11207 13515
rect 12526 13512 12532 13524
rect 11195 13484 12020 13512
rect 12487 13484 12532 13512
rect 11195 13481 11207 13484
rect 11149 13475 11207 13481
rect 5810 13404 5816 13456
rect 5868 13444 5874 13456
rect 7837 13447 7895 13453
rect 7837 13444 7849 13447
rect 5868 13416 7849 13444
rect 5868 13404 5874 13416
rect 7837 13413 7849 13416
rect 7883 13413 7895 13447
rect 7837 13407 7895 13413
rect 1670 13336 1676 13388
rect 1728 13376 1734 13388
rect 2225 13379 2283 13385
rect 2225 13376 2237 13379
rect 1728 13348 2237 13376
rect 1728 13336 1734 13348
rect 2225 13345 2237 13348
rect 2271 13345 2283 13379
rect 2225 13339 2283 13345
rect 4798 13336 4804 13388
rect 4856 13376 4862 13388
rect 4985 13379 5043 13385
rect 4985 13376 4997 13379
rect 4856 13348 4997 13376
rect 4856 13336 4862 13348
rect 4985 13345 4997 13348
rect 5031 13345 5043 13379
rect 4985 13339 5043 13345
rect 2133 13311 2191 13317
rect 2133 13277 2145 13311
rect 2179 13277 2191 13311
rect 2406 13308 2412 13320
rect 2367 13280 2412 13308
rect 2133 13271 2191 13277
rect 2148 13240 2176 13271
rect 2406 13268 2412 13280
rect 2464 13268 2470 13320
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13308 2559 13311
rect 3142 13308 3148 13320
rect 2547 13280 3148 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 5000 13308 5028 13339
rect 5261 13311 5319 13317
rect 5261 13308 5273 13311
rect 5000 13280 5273 13308
rect 5261 13277 5273 13280
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 5350 13268 5356 13320
rect 5408 13308 5414 13320
rect 6917 13311 6975 13317
rect 5408 13280 5453 13308
rect 5408 13268 5414 13280
rect 6917 13277 6929 13311
rect 6963 13308 6975 13311
rect 7006 13308 7012 13320
rect 6963 13280 7012 13308
rect 6963 13277 6975 13280
rect 6917 13271 6975 13277
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 8019 13317 8047 13472
rect 8297 13379 8355 13385
rect 8297 13345 8309 13379
rect 8343 13376 8355 13379
rect 9585 13379 9643 13385
rect 8343 13348 9260 13376
rect 8343 13345 8355 13348
rect 8297 13339 8355 13345
rect 9232 13320 9260 13348
rect 9585 13345 9597 13379
rect 9631 13376 9643 13379
rect 11882 13376 11888 13388
rect 9631 13348 11888 13376
rect 9631 13345 9643 13348
rect 9585 13339 9643 13345
rect 8019 13311 8079 13317
rect 8019 13280 8033 13311
rect 8021 13277 8033 13280
rect 8067 13277 8079 13311
rect 8021 13271 8079 13277
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13286 8171 13311
rect 8389 13311 8447 13317
rect 8159 13277 8248 13286
rect 8113 13271 8248 13277
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 8435 13280 9137 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 9125 13277 9137 13280
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 2774 13240 2780 13252
rect 2148 13212 2780 13240
rect 2774 13200 2780 13212
rect 2832 13200 2838 13252
rect 4706 13200 4712 13252
rect 4764 13240 4770 13252
rect 4893 13243 4951 13249
rect 4893 13240 4905 13243
rect 4764 13212 4905 13240
rect 4764 13200 4770 13212
rect 4893 13209 4905 13212
rect 4939 13240 4951 13243
rect 5368 13240 5396 13268
rect 8128 13258 8248 13271
rect 4939 13212 5396 13240
rect 8220 13240 8248 13258
rect 8938 13240 8944 13252
rect 8220 13212 8944 13240
rect 4939 13209 4951 13212
rect 4893 13203 4951 13209
rect 8938 13200 8944 13212
rect 8996 13200 9002 13252
rect 9140 13240 9168 13271
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 9493 13311 9551 13317
rect 9493 13308 9505 13311
rect 9272 13280 9505 13308
rect 9272 13268 9278 13280
rect 9493 13277 9505 13280
rect 9539 13277 9551 13311
rect 9493 13271 9551 13277
rect 9600 13240 9628 13339
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 11992 13385 12020 13484
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 13357 13515 13415 13521
rect 13357 13481 13369 13515
rect 13403 13512 13415 13515
rect 13538 13512 13544 13524
rect 13403 13484 13544 13512
rect 13403 13481 13415 13484
rect 13357 13475 13415 13481
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 14734 13512 14740 13524
rect 14695 13484 14740 13512
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 14182 13404 14188 13456
rect 14240 13444 14246 13456
rect 14277 13447 14335 13453
rect 14277 13444 14289 13447
rect 14240 13416 14289 13444
rect 14240 13404 14246 13416
rect 14277 13413 14289 13416
rect 14323 13413 14335 13447
rect 14277 13407 14335 13413
rect 11977 13379 12035 13385
rect 11977 13345 11989 13379
rect 12023 13345 12035 13379
rect 11977 13339 12035 13345
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 10505 13311 10563 13317
rect 10505 13308 10517 13311
rect 10284 13280 10517 13308
rect 10284 13268 10290 13280
rect 10505 13277 10517 13280
rect 10551 13277 10563 13311
rect 10505 13271 10563 13277
rect 10594 13268 10600 13320
rect 10652 13308 10658 13320
rect 10870 13308 10876 13320
rect 10652 13280 10876 13308
rect 10652 13268 10658 13280
rect 10870 13268 10876 13280
rect 10928 13308 10934 13320
rect 11179 13311 11237 13317
rect 11179 13308 11191 13311
rect 10928 13280 11191 13308
rect 10928 13268 10934 13280
rect 11179 13277 11191 13280
rect 11225 13277 11237 13311
rect 11179 13271 11237 13277
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 11992 13308 12020 13339
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 12345 13379 12403 13385
rect 12345 13376 12357 13379
rect 12216 13348 12357 13376
rect 12216 13336 12222 13348
rect 12345 13345 12357 13348
rect 12391 13345 12403 13379
rect 12345 13339 12403 13345
rect 12253 13311 12311 13317
rect 12253 13308 12265 13311
rect 11388 13280 11433 13308
rect 11992 13280 12265 13308
rect 11388 13268 11394 13280
rect 12253 13277 12265 13280
rect 12299 13277 12311 13311
rect 12434 13308 12440 13320
rect 12253 13271 12311 13277
rect 9140 13212 9628 13240
rect 10042 13200 10048 13252
rect 10100 13240 10106 13252
rect 11882 13240 11888 13252
rect 10100 13212 10456 13240
rect 11843 13212 11888 13240
rect 10100 13200 10106 13212
rect 10318 13172 10324 13184
rect 10279 13144 10324 13172
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 10428 13172 10456 13212
rect 11882 13200 11888 13212
rect 11940 13240 11946 13252
rect 12158 13240 12164 13252
rect 11940 13212 12164 13240
rect 11940 13200 11946 13212
rect 12158 13200 12164 13212
rect 12216 13200 12222 13252
rect 12268 13240 12296 13271
rect 12406 13268 12440 13308
rect 12492 13268 12498 13320
rect 12894 13268 12900 13320
rect 12952 13308 12958 13320
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 12952 13280 13185 13308
rect 12952 13268 12958 13280
rect 13173 13277 13185 13280
rect 13219 13308 13231 13311
rect 13630 13308 13636 13320
rect 13219 13280 13636 13308
rect 13219 13277 13231 13280
rect 13173 13271 13231 13277
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 14090 13268 14096 13320
rect 14148 13308 14154 13320
rect 14185 13311 14243 13317
rect 14185 13308 14197 13311
rect 14148 13280 14197 13308
rect 14148 13268 14154 13280
rect 14185 13277 14197 13280
rect 14231 13277 14243 13311
rect 14458 13308 14464 13320
rect 14419 13280 14464 13308
rect 14185 13271 14243 13277
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13308 14611 13311
rect 14642 13308 14648 13320
rect 14599 13280 14648 13308
rect 14599 13277 14611 13280
rect 14553 13271 14611 13277
rect 14642 13268 14648 13280
rect 14700 13268 14706 13320
rect 12406 13240 12434 13268
rect 12268 13212 12434 13240
rect 12989 13243 13047 13249
rect 12989 13209 13001 13243
rect 13035 13209 13047 13243
rect 12989 13203 13047 13209
rect 13004 13172 13032 13203
rect 10428 13144 13032 13172
rect 1104 13082 15732 13104
rect 1104 13030 5858 13082
rect 5910 13030 5922 13082
rect 5974 13030 5986 13082
rect 6038 13030 6050 13082
rect 6102 13030 10734 13082
rect 10786 13030 10798 13082
rect 10850 13030 10862 13082
rect 10914 13030 10926 13082
rect 10978 13030 15732 13082
rect 1104 13008 15732 13030
rect 2225 12971 2283 12977
rect 2225 12937 2237 12971
rect 2271 12968 2283 12971
rect 2406 12968 2412 12980
rect 2271 12940 2412 12968
rect 2271 12937 2283 12940
rect 2225 12931 2283 12937
rect 2406 12928 2412 12940
rect 2464 12928 2470 12980
rect 3513 12971 3571 12977
rect 3513 12937 3525 12971
rect 3559 12968 3571 12971
rect 5074 12968 5080 12980
rect 3559 12940 5080 12968
rect 3559 12937 3571 12940
rect 3513 12931 3571 12937
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 5718 12968 5724 12980
rect 5679 12940 5724 12968
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 11977 12971 12035 12977
rect 11977 12937 11989 12971
rect 12023 12968 12035 12971
rect 12023 12940 12434 12968
rect 12023 12937 12035 12940
rect 11977 12931 12035 12937
rect 1581 12903 1639 12909
rect 1581 12869 1593 12903
rect 1627 12900 1639 12903
rect 2961 12903 3019 12909
rect 1627 12872 2084 12900
rect 1627 12869 1639 12872
rect 1581 12863 1639 12869
rect 1949 12835 2007 12841
rect 1949 12832 1961 12835
rect 1688 12804 1961 12832
rect 1688 12776 1716 12804
rect 1949 12801 1961 12804
rect 1995 12801 2007 12835
rect 1949 12795 2007 12801
rect 1670 12724 1676 12776
rect 1728 12764 1734 12776
rect 2056 12773 2084 12872
rect 2961 12869 2973 12903
rect 3007 12900 3019 12903
rect 3007 12872 3280 12900
rect 3007 12869 3019 12872
rect 2961 12863 3019 12869
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 3050 12832 3056 12844
rect 2915 12804 3056 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 3252 12841 3280 12872
rect 8018 12860 8024 12912
rect 8076 12900 8082 12912
rect 10042 12900 10048 12912
rect 8076 12872 10048 12900
rect 8076 12860 8082 12872
rect 10042 12860 10048 12872
rect 10100 12860 10106 12912
rect 10244 12872 10456 12900
rect 3237 12835 3295 12841
rect 3237 12801 3249 12835
rect 3283 12832 3295 12835
rect 4249 12835 4307 12841
rect 3283 12804 4016 12832
rect 3283 12801 3295 12804
rect 3237 12795 3295 12801
rect 2041 12767 2099 12773
rect 1728 12736 1773 12764
rect 1728 12724 1734 12736
rect 2041 12733 2053 12767
rect 2087 12764 2099 12767
rect 2774 12764 2780 12776
rect 2087 12736 2780 12764
rect 2087 12733 2099 12736
rect 2041 12727 2099 12733
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 3068 12764 3096 12792
rect 3329 12767 3387 12773
rect 3329 12764 3341 12767
rect 3068 12736 3341 12764
rect 3329 12733 3341 12736
rect 3375 12733 3387 12767
rect 3329 12727 3387 12733
rect 3988 12637 4016 12804
rect 4249 12801 4261 12835
rect 4295 12801 4307 12835
rect 4249 12795 4307 12801
rect 4157 12767 4215 12773
rect 4157 12733 4169 12767
rect 4203 12733 4215 12767
rect 4264 12764 4292 12795
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5776 12804 5825 12832
rect 5776 12792 5782 12804
rect 5813 12801 5825 12804
rect 5859 12832 5871 12835
rect 6178 12832 6184 12844
rect 5859 12804 6184 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 6546 12832 6552 12844
rect 6507 12804 6552 12832
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7466 12832 7472 12844
rect 7156 12804 7472 12832
rect 7156 12792 7162 12804
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 9214 12832 9220 12844
rect 9175 12804 9220 12832
rect 9214 12792 9220 12804
rect 9272 12792 9278 12844
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12832 9459 12835
rect 9766 12832 9772 12844
rect 9447 12804 9772 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 9950 12832 9956 12844
rect 9911 12804 9956 12832
rect 9950 12792 9956 12804
rect 10008 12792 10014 12844
rect 10244 12841 10272 12872
rect 10229 12835 10287 12841
rect 10229 12801 10241 12835
rect 10275 12801 10287 12835
rect 10229 12795 10287 12801
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12801 10379 12835
rect 10428 12832 10456 12872
rect 10502 12860 10508 12912
rect 10560 12900 10566 12912
rect 12406 12900 12434 12940
rect 14458 12928 14464 12980
rect 14516 12968 14522 12980
rect 14737 12971 14795 12977
rect 14737 12968 14749 12971
rect 14516 12940 14749 12968
rect 14516 12928 14522 12940
rect 14737 12937 14749 12940
rect 14783 12937 14795 12971
rect 14737 12931 14795 12937
rect 13722 12900 13728 12912
rect 10560 12872 12296 12900
rect 12406 12872 13728 12900
rect 10560 12860 10566 12872
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 10428 12804 11529 12832
rect 10321 12795 10379 12801
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 4430 12764 4436 12776
rect 4264 12736 4436 12764
rect 4157 12727 4215 12733
rect 4172 12696 4200 12727
rect 4430 12724 4436 12736
rect 4488 12764 4494 12776
rect 4525 12767 4583 12773
rect 4525 12764 4537 12767
rect 4488 12736 4537 12764
rect 4488 12724 4494 12736
rect 4525 12733 4537 12736
rect 4571 12733 4583 12767
rect 4525 12727 4583 12733
rect 4617 12767 4675 12773
rect 4617 12733 4629 12767
rect 4663 12764 4675 12767
rect 7006 12764 7012 12776
rect 4663 12736 7012 12764
rect 4663 12733 4675 12736
rect 4617 12727 4675 12733
rect 4338 12696 4344 12708
rect 4172 12668 4344 12696
rect 4338 12656 4344 12668
rect 4396 12696 4402 12708
rect 4632 12696 4660 12727
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12764 7803 12767
rect 9490 12764 9496 12776
rect 7791 12736 9496 12764
rect 7791 12733 7803 12736
rect 7745 12727 7803 12733
rect 9490 12724 9496 12736
rect 9548 12724 9554 12776
rect 4396 12668 4660 12696
rect 4396 12656 4402 12668
rect 8662 12656 8668 12708
rect 8720 12696 8726 12708
rect 10244 12696 10272 12795
rect 10336 12764 10364 12795
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 11793 12835 11851 12841
rect 11793 12832 11805 12835
rect 11756 12804 11805 12832
rect 11756 12792 11762 12804
rect 11793 12801 11805 12804
rect 11839 12801 11851 12835
rect 11793 12795 11851 12801
rect 11974 12792 11980 12844
rect 12032 12832 12038 12844
rect 12158 12832 12164 12844
rect 12032 12804 12164 12832
rect 12032 12792 12038 12804
rect 12158 12792 12164 12804
rect 12216 12792 12222 12844
rect 12268 12832 12296 12872
rect 13188 12841 13216 12872
rect 13722 12860 13728 12872
rect 13780 12860 13786 12912
rect 12437 12835 12495 12841
rect 12437 12832 12449 12835
rect 12268 12804 12449 12832
rect 12437 12801 12449 12804
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12801 13231 12835
rect 13173 12795 13231 12801
rect 14461 12835 14519 12841
rect 14461 12801 14473 12835
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 10686 12764 10692 12776
rect 10336 12736 10692 12764
rect 10686 12724 10692 12736
rect 10744 12764 10750 12776
rect 11609 12767 11667 12773
rect 11609 12764 11621 12767
rect 10744 12736 11621 12764
rect 10744 12724 10750 12736
rect 11609 12733 11621 12736
rect 11655 12733 11667 12767
rect 11609 12727 11667 12733
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 14090 12764 14096 12776
rect 13679 12736 14096 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 14090 12724 14096 12736
rect 14148 12724 14154 12776
rect 14182 12724 14188 12776
rect 14240 12764 14246 12776
rect 14476 12764 14504 12795
rect 14240 12736 14504 12764
rect 14553 12767 14611 12773
rect 14240 12724 14246 12736
rect 14553 12733 14565 12767
rect 14599 12733 14611 12767
rect 14553 12727 14611 12733
rect 8720 12668 10272 12696
rect 10505 12699 10563 12705
rect 8720 12656 8726 12668
rect 10505 12665 10517 12699
rect 10551 12696 10563 12699
rect 14108 12696 14136 12724
rect 14568 12696 14596 12727
rect 10551 12668 13308 12696
rect 14108 12668 14596 12696
rect 10551 12665 10563 12668
rect 10505 12659 10563 12665
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 4062 12628 4068 12640
rect 4019 12600 4068 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 6641 12631 6699 12637
rect 6641 12628 6653 12631
rect 6604 12600 6653 12628
rect 6604 12588 6610 12600
rect 6641 12597 6653 12600
rect 6687 12597 6699 12631
rect 6641 12591 6699 12597
rect 8846 12588 8852 12640
rect 8904 12628 8910 12640
rect 9033 12631 9091 12637
rect 9033 12628 9045 12631
rect 8904 12600 9045 12628
rect 8904 12588 8910 12600
rect 9033 12597 9045 12600
rect 9079 12597 9091 12631
rect 9033 12591 9091 12597
rect 10045 12631 10103 12637
rect 10045 12597 10057 12631
rect 10091 12628 10103 12631
rect 10134 12628 10140 12640
rect 10091 12600 10140 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 11790 12628 11796 12640
rect 11751 12600 11796 12628
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 13280 12637 13308 12668
rect 12621 12631 12679 12637
rect 12621 12628 12633 12631
rect 12492 12600 12633 12628
rect 12492 12588 12498 12600
rect 12621 12597 12633 12600
rect 12667 12597 12679 12631
rect 12621 12591 12679 12597
rect 13265 12631 13323 12637
rect 13265 12597 13277 12631
rect 13311 12597 13323 12631
rect 13265 12591 13323 12597
rect 1104 12538 15732 12560
rect 1104 12486 3420 12538
rect 3472 12486 3484 12538
rect 3536 12486 3548 12538
rect 3600 12486 3612 12538
rect 3664 12486 8296 12538
rect 8348 12486 8360 12538
rect 8412 12486 8424 12538
rect 8476 12486 8488 12538
rect 8540 12486 13172 12538
rect 13224 12486 13236 12538
rect 13288 12486 13300 12538
rect 13352 12486 13364 12538
rect 13416 12486 15732 12538
rect 1104 12464 15732 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 2832 12396 3801 12424
rect 2832 12384 2838 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 5350 12424 5356 12436
rect 5311 12396 5356 12424
rect 3789 12387 3847 12393
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 7190 12424 7196 12436
rect 7151 12396 7196 12424
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 7650 12424 7656 12436
rect 7563 12396 7656 12424
rect 7650 12384 7656 12396
rect 7708 12424 7714 12436
rect 8018 12424 8024 12436
rect 7708 12396 8024 12424
rect 7708 12384 7714 12396
rect 8018 12384 8024 12396
rect 8076 12384 8082 12436
rect 8205 12427 8263 12433
rect 8205 12393 8217 12427
rect 8251 12424 8263 12427
rect 8662 12424 8668 12436
rect 8251 12396 8668 12424
rect 8251 12393 8263 12396
rect 8205 12387 8263 12393
rect 8312 12368 8340 12396
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 9214 12424 9220 12436
rect 9175 12396 9220 12424
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 9950 12424 9956 12436
rect 9692 12396 9956 12424
rect 8294 12316 8300 12368
rect 8352 12316 8358 12368
rect 4249 12291 4307 12297
rect 4249 12257 4261 12291
rect 4295 12288 4307 12291
rect 4430 12288 4436 12300
rect 4295 12260 4436 12288
rect 4295 12257 4307 12260
rect 4249 12251 4307 12257
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 7098 12248 7104 12300
rect 7156 12288 7162 12300
rect 7156 12260 8432 12288
rect 7156 12248 7162 12260
rect 3050 12180 3056 12232
rect 3108 12220 3114 12232
rect 3970 12220 3976 12232
rect 3108 12192 3976 12220
rect 3108 12180 3114 12192
rect 3970 12180 3976 12192
rect 4028 12180 4034 12232
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4338 12220 4344 12232
rect 4120 12192 4165 12220
rect 4299 12192 4344 12220
rect 4120 12180 4126 12192
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 5552 12152 5580 12183
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 5905 12223 5963 12229
rect 5905 12220 5917 12223
rect 5684 12192 5917 12220
rect 5684 12180 5690 12192
rect 5905 12189 5917 12192
rect 5951 12189 5963 12223
rect 6546 12220 6552 12232
rect 6507 12192 6552 12220
rect 5905 12183 5963 12189
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 7374 12220 7380 12232
rect 7335 12192 7380 12220
rect 7374 12180 7380 12192
rect 7432 12180 7438 12232
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 7745 12223 7803 12229
rect 7524 12192 7569 12220
rect 7524 12180 7530 12192
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 8294 12220 8300 12232
rect 7791 12192 8300 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8404 12229 8432 12260
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 9692 12297 9720 12396
rect 9950 12384 9956 12396
rect 10008 12424 10014 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 10008 12396 10241 12424
rect 10008 12384 10014 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 11882 12424 11888 12436
rect 11843 12396 11888 12424
rect 10229 12387 10287 12393
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 13541 12427 13599 12433
rect 13541 12393 13553 12427
rect 13587 12424 13599 12427
rect 14182 12424 14188 12436
rect 13587 12396 14188 12424
rect 13587 12393 13599 12396
rect 13541 12387 13599 12393
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 14737 12427 14795 12433
rect 14737 12393 14749 12427
rect 14783 12424 14795 12427
rect 14826 12424 14832 12436
rect 14783 12396 14832 12424
rect 14783 12393 14795 12396
rect 14737 12387 14795 12393
rect 14826 12384 14832 12396
rect 14884 12384 14890 12436
rect 9766 12316 9772 12368
rect 9824 12356 9830 12368
rect 10689 12359 10747 12365
rect 10689 12356 10701 12359
rect 9824 12328 10701 12356
rect 9824 12316 9830 12328
rect 10689 12325 10701 12328
rect 10735 12356 10747 12359
rect 14642 12356 14648 12368
rect 10735 12328 14648 12356
rect 10735 12325 10747 12328
rect 10689 12319 10747 12325
rect 9677 12291 9735 12297
rect 9677 12288 9689 12291
rect 8536 12260 9689 12288
rect 8536 12248 8542 12260
rect 9677 12257 9689 12260
rect 9723 12257 9735 12291
rect 9677 12251 9735 12257
rect 9950 12248 9956 12300
rect 10008 12288 10014 12300
rect 10321 12291 10379 12297
rect 10321 12288 10333 12291
rect 10008 12260 10333 12288
rect 10008 12248 10014 12260
rect 10321 12257 10333 12260
rect 10367 12288 10379 12291
rect 12894 12288 12900 12300
rect 10367 12260 12900 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 12894 12248 12900 12260
rect 12952 12288 12958 12300
rect 14476 12297 14504 12328
rect 14642 12316 14648 12328
rect 14700 12316 14706 12368
rect 14461 12291 14519 12297
rect 12952 12260 13400 12288
rect 12952 12248 12958 12260
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 9306 12220 9312 12232
rect 9088 12192 9312 12220
rect 9088 12180 9094 12192
rect 9306 12180 9312 12192
rect 9364 12220 9370 12232
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 9364 12192 9413 12220
rect 9364 12180 9370 12192
rect 9401 12189 9413 12192
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12189 9551 12223
rect 9766 12220 9772 12232
rect 9679 12192 9772 12220
rect 9493 12183 9551 12189
rect 5997 12155 6055 12161
rect 5997 12152 6009 12155
rect 5552 12124 6009 12152
rect 5997 12121 6009 12124
rect 6043 12152 6055 12155
rect 6178 12152 6184 12164
rect 6043 12124 6184 12152
rect 6043 12121 6055 12124
rect 5997 12115 6055 12121
rect 6178 12112 6184 12124
rect 6236 12112 6242 12164
rect 9508 12152 9536 12183
rect 9766 12180 9772 12192
rect 9824 12220 9830 12232
rect 10505 12223 10563 12229
rect 10505 12220 10517 12223
rect 9824 12192 10517 12220
rect 9824 12180 9830 12192
rect 10505 12189 10517 12192
rect 10551 12220 10563 12223
rect 10686 12220 10692 12232
rect 10551 12192 10692 12220
rect 10551 12189 10563 12192
rect 10505 12183 10563 12189
rect 10686 12180 10692 12192
rect 10744 12220 10750 12232
rect 11146 12220 11152 12232
rect 10744 12192 11152 12220
rect 10744 12180 10750 12192
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 11698 12220 11704 12232
rect 11659 12192 11704 12220
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 13372 12229 13400 12260
rect 14461 12257 14473 12291
rect 14507 12288 14519 12291
rect 15013 12291 15071 12297
rect 15013 12288 15025 12291
rect 14507 12260 15025 12288
rect 14507 12257 14519 12260
rect 14461 12251 14519 12257
rect 15013 12257 15025 12260
rect 15059 12257 15071 12291
rect 15013 12251 15071 12257
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 12452 12192 13185 12220
rect 12452 12164 12480 12192
rect 13173 12189 13185 12192
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12189 13415 12223
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 13357 12183 13415 12189
rect 14568 12192 14841 12220
rect 10229 12155 10287 12161
rect 10229 12152 10241 12155
rect 9508 12124 10241 12152
rect 10229 12121 10241 12124
rect 10275 12121 10287 12155
rect 10229 12115 10287 12121
rect 6733 12087 6791 12093
rect 6733 12053 6745 12087
rect 6779 12084 6791 12087
rect 7374 12084 7380 12096
rect 6779 12056 7380 12084
rect 6779 12053 6791 12056
rect 6733 12047 6791 12053
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 10134 12044 10140 12096
rect 10192 12084 10198 12096
rect 10244 12084 10272 12115
rect 11422 12112 11428 12164
rect 11480 12152 11486 12164
rect 11517 12155 11575 12161
rect 11517 12152 11529 12155
rect 11480 12124 11529 12152
rect 11480 12112 11486 12124
rect 11517 12121 11529 12124
rect 11563 12152 11575 12155
rect 12345 12155 12403 12161
rect 12345 12152 12357 12155
rect 11563 12124 12357 12152
rect 11563 12121 11575 12124
rect 11517 12115 11575 12121
rect 12345 12121 12357 12124
rect 12391 12152 12403 12155
rect 12434 12152 12440 12164
rect 12391 12124 12440 12152
rect 12391 12121 12403 12124
rect 12345 12115 12403 12121
rect 12434 12112 12440 12124
rect 12492 12112 12498 12164
rect 12529 12155 12587 12161
rect 12529 12121 12541 12155
rect 12575 12121 12587 12155
rect 12529 12115 12587 12121
rect 11790 12084 11796 12096
rect 10192 12056 11796 12084
rect 10192 12044 10198 12056
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 11974 12044 11980 12096
rect 12032 12084 12038 12096
rect 12544 12084 12572 12115
rect 12032 12056 12572 12084
rect 12713 12087 12771 12093
rect 12032 12044 12038 12056
rect 12713 12053 12725 12087
rect 12759 12084 12771 12087
rect 12894 12084 12900 12096
rect 12759 12056 12900 12084
rect 12759 12053 12771 12056
rect 12713 12047 12771 12053
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 14568 12093 14596 12192
rect 14829 12189 14841 12192
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 14553 12087 14611 12093
rect 14553 12084 14565 12087
rect 14516 12056 14565 12084
rect 14516 12044 14522 12056
rect 14553 12053 14565 12056
rect 14599 12053 14611 12087
rect 14553 12047 14611 12053
rect 1104 11994 15732 12016
rect 1104 11942 5858 11994
rect 5910 11942 5922 11994
rect 5974 11942 5986 11994
rect 6038 11942 6050 11994
rect 6102 11942 10734 11994
rect 10786 11942 10798 11994
rect 10850 11942 10862 11994
rect 10914 11942 10926 11994
rect 10978 11942 15732 11994
rect 1104 11920 15732 11942
rect 1670 11880 1676 11892
rect 1631 11852 1676 11880
rect 1670 11840 1676 11852
rect 1728 11840 1734 11892
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 7193 11883 7251 11889
rect 7193 11880 7205 11883
rect 7064 11852 7205 11880
rect 7064 11840 7070 11852
rect 7193 11849 7205 11852
rect 7239 11849 7251 11883
rect 8018 11880 8024 11892
rect 7931 11852 8024 11880
rect 7193 11843 7251 11849
rect 8018 11840 8024 11852
rect 8076 11880 8082 11892
rect 8478 11880 8484 11892
rect 8076 11852 8484 11880
rect 8076 11840 8082 11852
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 9950 11880 9956 11892
rect 9232 11852 9956 11880
rect 4341 11815 4399 11821
rect 4341 11781 4353 11815
rect 4387 11812 4399 11815
rect 6730 11812 6736 11824
rect 4387 11784 5488 11812
rect 6691 11784 6736 11812
rect 4387 11781 4399 11784
rect 4341 11775 4399 11781
rect 1946 11744 1952 11756
rect 1907 11716 1952 11744
rect 1946 11704 1952 11716
rect 2004 11744 2010 11756
rect 2225 11747 2283 11753
rect 2225 11744 2237 11747
rect 2004 11716 2237 11744
rect 2004 11704 2010 11716
rect 2225 11713 2237 11716
rect 2271 11713 2283 11747
rect 2225 11707 2283 11713
rect 3234 11704 3240 11756
rect 3292 11744 3298 11756
rect 3605 11747 3663 11753
rect 3605 11744 3617 11747
rect 3292 11716 3617 11744
rect 3292 11704 3298 11716
rect 3605 11713 3617 11716
rect 3651 11713 3663 11747
rect 3786 11744 3792 11756
rect 3747 11716 3792 11744
rect 3605 11707 3663 11713
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 3881 11747 3939 11753
rect 3881 11713 3893 11747
rect 3927 11744 3939 11747
rect 4154 11744 4160 11756
rect 3927 11716 4160 11744
rect 3927 11713 3939 11716
rect 3881 11707 3939 11713
rect 4154 11704 4160 11716
rect 4212 11704 4218 11756
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11713 4583 11747
rect 4525 11707 4583 11713
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 5258 11744 5264 11756
rect 4755 11716 5264 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 1857 11679 1915 11685
rect 1857 11645 1869 11679
rect 1903 11676 1915 11679
rect 2317 11679 2375 11685
rect 2317 11676 2329 11679
rect 1903 11648 2329 11676
rect 1903 11645 1915 11648
rect 1857 11639 1915 11645
rect 2317 11645 2329 11648
rect 2363 11676 2375 11679
rect 2958 11676 2964 11688
rect 2363 11648 2964 11676
rect 2363 11645 2375 11648
rect 2317 11639 2375 11645
rect 2958 11636 2964 11648
rect 3016 11636 3022 11688
rect 4540 11676 4568 11707
rect 5258 11704 5264 11716
rect 5316 11744 5322 11756
rect 5353 11747 5411 11753
rect 5353 11744 5365 11747
rect 5316 11716 5365 11744
rect 5316 11704 5322 11716
rect 5353 11713 5365 11716
rect 5399 11713 5411 11747
rect 5460 11744 5488 11784
rect 6730 11772 6736 11784
rect 6788 11772 6794 11824
rect 8849 11815 8907 11821
rect 8849 11812 8861 11815
rect 6840 11784 8861 11812
rect 5626 11753 5632 11756
rect 5582 11747 5632 11753
rect 5582 11744 5594 11747
rect 5460 11716 5594 11744
rect 5353 11707 5411 11713
rect 5582 11713 5594 11716
rect 5628 11713 5632 11747
rect 5582 11707 5632 11713
rect 5626 11704 5632 11707
rect 5684 11704 5690 11756
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6178 11744 6184 11756
rect 5859 11716 6184 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 6178 11704 6184 11716
rect 6236 11744 6242 11756
rect 6840 11744 6868 11784
rect 8849 11781 8861 11784
rect 8895 11781 8907 11815
rect 8849 11775 8907 11781
rect 7006 11744 7012 11756
rect 6236 11716 6868 11744
rect 6967 11716 7012 11744
rect 6236 11704 6242 11716
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 7374 11704 7380 11756
rect 7432 11744 7438 11756
rect 7837 11747 7895 11753
rect 7837 11744 7849 11747
rect 7432 11716 7849 11744
rect 7432 11704 7438 11716
rect 7837 11713 7849 11716
rect 7883 11713 7895 11747
rect 7837 11707 7895 11713
rect 6454 11676 6460 11688
rect 4540 11648 6460 11676
rect 6454 11636 6460 11648
rect 6512 11636 6518 11688
rect 6546 11636 6552 11688
rect 6604 11676 6610 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6604 11648 6837 11676
rect 6604 11636 6610 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 3050 11568 3056 11620
rect 3108 11608 3114 11620
rect 5169 11611 5227 11617
rect 5169 11608 5181 11611
rect 3108 11580 5181 11608
rect 3108 11568 3114 11580
rect 5169 11577 5181 11580
rect 5215 11577 5227 11611
rect 7742 11608 7748 11620
rect 5169 11571 5227 11577
rect 6840 11580 7748 11608
rect 3605 11543 3663 11549
rect 3605 11509 3617 11543
rect 3651 11540 3663 11543
rect 3878 11540 3884 11552
rect 3651 11512 3884 11540
rect 3651 11509 3663 11512
rect 3605 11503 3663 11509
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 6840 11549 6868 11580
rect 7742 11568 7748 11580
rect 7800 11568 7806 11620
rect 7852 11608 7880 11707
rect 7926 11704 7932 11756
rect 7984 11744 7990 11756
rect 8110 11744 8116 11756
rect 7984 11716 8116 11744
rect 7984 11704 7990 11716
rect 8110 11704 8116 11716
rect 8168 11744 8174 11756
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 8168 11716 8493 11744
rect 8168 11704 8174 11716
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11744 8723 11747
rect 9232 11744 9260 11852
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 10134 11880 10140 11892
rect 10095 11852 10140 11880
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 10781 11883 10839 11889
rect 10781 11849 10793 11883
rect 10827 11880 10839 11883
rect 11146 11880 11152 11892
rect 10827 11852 11152 11880
rect 10827 11849 10839 11852
rect 10781 11843 10839 11849
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 11330 11840 11336 11892
rect 11388 11880 11394 11892
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 11388 11852 11529 11880
rect 11388 11840 11394 11852
rect 11517 11849 11529 11852
rect 11563 11849 11575 11883
rect 11517 11843 11575 11849
rect 9766 11812 9772 11824
rect 9508 11784 9772 11812
rect 9508 11753 9536 11784
rect 9766 11772 9772 11784
rect 9824 11772 9830 11824
rect 10686 11772 10692 11824
rect 10744 11812 10750 11824
rect 12894 11812 12900 11824
rect 10744 11784 11836 11812
rect 12855 11784 12900 11812
rect 10744 11772 10750 11784
rect 8711 11716 9260 11744
rect 9309 11747 9367 11753
rect 8711 11713 8723 11716
rect 8665 11707 8723 11713
rect 9309 11713 9321 11747
rect 9355 11713 9367 11747
rect 9309 11707 9367 11713
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 10321 11747 10379 11753
rect 10321 11713 10333 11747
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11744 11023 11747
rect 11514 11744 11520 11756
rect 11011 11716 11520 11744
rect 11011 11713 11023 11716
rect 10965 11707 11023 11713
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 9324 11676 9352 11707
rect 9088 11648 9352 11676
rect 10336 11676 10364 11707
rect 11514 11704 11520 11716
rect 11572 11744 11578 11756
rect 11808 11753 11836 11784
rect 12894 11772 12900 11784
rect 12952 11812 12958 11824
rect 12952 11784 13216 11812
rect 12952 11772 12958 11784
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11572 11716 11713 11744
rect 11572 11704 11578 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 13188 11753 13216 11784
rect 12069 11747 12127 11753
rect 12069 11744 12081 11747
rect 11940 11716 12081 11744
rect 11940 11704 11946 11716
rect 12069 11713 12081 11716
rect 12115 11713 12127 11747
rect 12069 11707 12127 11713
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 14090 11744 14096 11756
rect 14051 11716 14096 11744
rect 13173 11707 13231 11713
rect 14090 11704 14096 11716
rect 14148 11704 14154 11756
rect 14918 11744 14924 11756
rect 14879 11716 14924 11744
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 11146 11676 11152 11688
rect 10336 11648 11152 11676
rect 9088 11636 9094 11648
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 12802 11676 12808 11688
rect 12763 11648 12808 11676
rect 12802 11636 12808 11648
rect 12860 11676 12866 11688
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 12860 11648 13277 11676
rect 12860 11636 12866 11648
rect 13265 11645 13277 11648
rect 13311 11645 13323 11679
rect 13265 11639 13323 11645
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11676 14243 11679
rect 14826 11676 14832 11688
rect 14231 11648 14832 11676
rect 14231 11645 14243 11648
rect 14185 11639 14243 11645
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 11698 11608 11704 11620
rect 7852 11580 11704 11608
rect 11698 11568 11704 11580
rect 11756 11568 11762 11620
rect 13814 11568 13820 11620
rect 13872 11608 13878 11620
rect 14737 11611 14795 11617
rect 14737 11608 14749 11611
rect 13872 11580 14749 11608
rect 13872 11568 13878 11580
rect 14737 11577 14749 11580
rect 14783 11577 14795 11611
rect 14737 11571 14795 11577
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 7190 11500 7196 11552
rect 7248 11540 7254 11552
rect 8018 11540 8024 11552
rect 7248 11512 8024 11540
rect 7248 11500 7254 11512
rect 8018 11500 8024 11512
rect 8076 11500 8082 11552
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 9272 11512 9321 11540
rect 9272 11500 9278 11512
rect 9309 11509 9321 11512
rect 9355 11509 9367 11543
rect 9309 11503 9367 11509
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 10686 11540 10692 11552
rect 10376 11512 10692 11540
rect 10376 11500 10382 11512
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 11974 11540 11980 11552
rect 11935 11512 11980 11540
rect 11974 11500 11980 11512
rect 12032 11500 12038 11552
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 13449 11543 13507 11549
rect 13449 11540 13461 11543
rect 13044 11512 13461 11540
rect 13044 11500 13050 11512
rect 13449 11509 13461 11512
rect 13495 11509 13507 11543
rect 13449 11503 13507 11509
rect 1104 11450 15732 11472
rect 1104 11398 3420 11450
rect 3472 11398 3484 11450
rect 3536 11398 3548 11450
rect 3600 11398 3612 11450
rect 3664 11398 8296 11450
rect 8348 11398 8360 11450
rect 8412 11398 8424 11450
rect 8476 11398 8488 11450
rect 8540 11398 13172 11450
rect 13224 11398 13236 11450
rect 13288 11398 13300 11450
rect 13352 11398 13364 11450
rect 13416 11398 15732 11450
rect 1104 11376 15732 11398
rect 1489 11339 1547 11345
rect 1489 11305 1501 11339
rect 1535 11336 1547 11339
rect 1946 11336 1952 11348
rect 1535 11308 1952 11336
rect 1535 11305 1547 11308
rect 1489 11299 1547 11305
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 2685 11339 2743 11345
rect 2685 11305 2697 11339
rect 2731 11336 2743 11339
rect 3050 11336 3056 11348
rect 2731 11308 3056 11336
rect 2731 11305 2743 11308
rect 2685 11299 2743 11305
rect 3050 11296 3056 11308
rect 3108 11296 3114 11348
rect 3142 11296 3148 11348
rect 3200 11336 3206 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3200 11308 3801 11336
rect 3200 11296 3206 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 5258 11336 5264 11348
rect 5219 11308 5264 11336
rect 3789 11299 3847 11305
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 6512 11308 6561 11336
rect 6512 11296 6518 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 6549 11299 6607 11305
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 7156 11308 10548 11336
rect 7156 11296 7162 11308
rect 1964 11268 1992 11296
rect 1964 11240 2728 11268
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11200 1731 11203
rect 2038 11200 2044 11212
rect 1719 11172 2044 11200
rect 1719 11169 1731 11172
rect 1673 11163 1731 11169
rect 2038 11160 2044 11172
rect 2096 11200 2102 11212
rect 2133 11203 2191 11209
rect 2133 11200 2145 11203
rect 2096 11172 2145 11200
rect 2096 11160 2102 11172
rect 2133 11169 2145 11172
rect 2179 11169 2191 11203
rect 2133 11163 2191 11169
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11132 1823 11135
rect 2148 11132 2176 11163
rect 2593 11135 2651 11141
rect 2593 11132 2605 11135
rect 1811 11104 2084 11132
rect 2148 11104 2605 11132
rect 1811 11101 1823 11104
rect 1765 11095 1823 11101
rect 2056 11073 2084 11104
rect 2593 11101 2605 11104
rect 2639 11101 2651 11135
rect 2700 11132 2728 11240
rect 2809 11135 2867 11141
rect 2809 11132 2821 11135
rect 2700 11104 2821 11132
rect 2593 11095 2651 11101
rect 2809 11101 2821 11104
rect 2855 11101 2867 11135
rect 2958 11132 2964 11144
rect 2919 11104 2964 11132
rect 2809 11095 2867 11101
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 2041 11067 2099 11073
rect 2041 11033 2053 11067
rect 2087 11064 2099 11067
rect 3068 11064 3096 11296
rect 5626 11228 5632 11280
rect 5684 11268 5690 11280
rect 5813 11271 5871 11277
rect 5813 11268 5825 11271
rect 5684 11240 5825 11268
rect 5684 11228 5690 11240
rect 5813 11237 5825 11240
rect 5859 11237 5871 11271
rect 5813 11231 5871 11237
rect 7009 11271 7067 11277
rect 7009 11237 7021 11271
rect 7055 11268 7067 11271
rect 7466 11268 7472 11280
rect 7055 11240 7472 11268
rect 7055 11237 7067 11240
rect 7009 11231 7067 11237
rect 7466 11228 7472 11240
rect 7524 11268 7530 11280
rect 8110 11268 8116 11280
rect 7524 11240 8116 11268
rect 7524 11228 7530 11240
rect 8110 11228 8116 11240
rect 8168 11228 8174 11280
rect 9766 11228 9772 11280
rect 9824 11268 9830 11280
rect 10229 11271 10287 11277
rect 10229 11268 10241 11271
rect 9824 11240 10241 11268
rect 9824 11228 9830 11240
rect 10229 11237 10241 11240
rect 10275 11237 10287 11271
rect 10520 11268 10548 11308
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 10652 11308 10977 11336
rect 10652 11296 10658 11308
rect 10965 11305 10977 11308
rect 11011 11305 11023 11339
rect 10965 11299 11023 11305
rect 11149 11339 11207 11345
rect 11149 11305 11161 11339
rect 11195 11336 11207 11339
rect 11974 11336 11980 11348
rect 11195 11308 11980 11336
rect 11195 11305 11207 11308
rect 11149 11299 11207 11305
rect 11164 11268 11192 11299
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 12710 11336 12716 11348
rect 12671 11308 12716 11336
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 12894 11296 12900 11348
rect 12952 11336 12958 11348
rect 13173 11339 13231 11345
rect 13173 11336 13185 11339
rect 12952 11308 13185 11336
rect 12952 11296 12958 11308
rect 13173 11305 13185 11308
rect 13219 11305 13231 11339
rect 13173 11299 13231 11305
rect 13906 11296 13912 11348
rect 13964 11336 13970 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 13964 11308 14105 11336
rect 13964 11296 13970 11308
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 14093 11299 14151 11305
rect 14734 11296 14740 11348
rect 14792 11296 14798 11348
rect 10520 11240 11192 11268
rect 12253 11271 12311 11277
rect 10229 11231 10287 11237
rect 12253 11237 12265 11271
rect 12299 11268 12311 11271
rect 12802 11268 12808 11280
rect 12299 11240 12808 11268
rect 12299 11237 12311 11240
rect 12253 11231 12311 11237
rect 12802 11228 12808 11240
rect 12860 11268 12866 11280
rect 12860 11240 13032 11268
rect 12860 11228 12866 11240
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 3988 11172 4445 11200
rect 3602 11092 3608 11144
rect 3660 11132 3666 11144
rect 3786 11132 3792 11144
rect 3660 11104 3792 11132
rect 3660 11092 3666 11104
rect 3786 11092 3792 11104
rect 3844 11132 3850 11144
rect 3988 11141 4016 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 7374 11200 7380 11212
rect 4433 11163 4491 11169
rect 6748 11172 7380 11200
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3844 11104 3985 11132
rect 3844 11092 3850 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11132 4123 11135
rect 4154 11132 4160 11144
rect 4111 11104 4160 11132
rect 4111 11101 4123 11104
rect 4065 11095 4123 11101
rect 4154 11092 4160 11104
rect 4212 11132 4218 11144
rect 5629 11135 5687 11141
rect 4212 11104 4384 11132
rect 4212 11092 4218 11104
rect 2087 11036 3096 11064
rect 2087 11033 2099 11036
rect 2041 11027 2099 11033
rect 3142 11024 3148 11076
rect 3200 11064 3206 11076
rect 4356 11073 4384 11104
rect 5629 11101 5641 11135
rect 5675 11132 5687 11135
rect 5718 11132 5724 11144
rect 5675 11104 5724 11132
rect 5675 11101 5687 11104
rect 5629 11095 5687 11101
rect 5718 11092 5724 11104
rect 5776 11092 5782 11144
rect 6748 11141 6776 11172
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 7561 11203 7619 11209
rect 7561 11169 7573 11203
rect 7607 11200 7619 11203
rect 8662 11200 8668 11212
rect 7607 11172 8668 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11101 6883 11135
rect 6825 11095 6883 11101
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 7576 11132 7604 11163
rect 8662 11160 8668 11172
rect 8720 11160 8726 11212
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11200 11391 11203
rect 11514 11200 11520 11212
rect 11379 11172 11520 11200
rect 11379 11169 11391 11172
rect 11333 11163 11391 11169
rect 11514 11160 11520 11172
rect 11572 11160 11578 11212
rect 12342 11200 12348 11212
rect 11716 11172 12348 11200
rect 7834 11132 7840 11144
rect 7147 11104 7604 11132
rect 7795 11104 7840 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 4341 11067 4399 11073
rect 3200 11036 3245 11064
rect 3200 11024 3206 11036
rect 4341 11033 4353 11067
rect 4387 11064 4399 11067
rect 4982 11064 4988 11076
rect 4387 11036 4988 11064
rect 4387 11033 4399 11036
rect 4341 11027 4399 11033
rect 4982 11024 4988 11036
rect 5040 11024 5046 11076
rect 5534 11064 5540 11076
rect 5447 11036 5540 11064
rect 5534 11024 5540 11036
rect 5592 11064 5598 11076
rect 6270 11064 6276 11076
rect 5592 11036 6276 11064
rect 5592 11024 5598 11036
rect 6270 11024 6276 11036
rect 6328 11024 6334 11076
rect 6840 11064 6868 11095
rect 7834 11092 7840 11104
rect 7892 11092 7898 11144
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8904 11104 9137 11132
rect 8904 11092 8910 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 11146 11132 11152 11144
rect 11107 11104 11152 11132
rect 9125 11095 9183 11101
rect 11146 11092 11152 11104
rect 11204 11132 11210 11144
rect 11716 11132 11744 11172
rect 12342 11160 12348 11172
rect 12400 11160 12406 11212
rect 13004 11200 13032 11240
rect 13078 11228 13084 11280
rect 13136 11268 13142 11280
rect 13630 11268 13636 11280
rect 13136 11240 13636 11268
rect 13136 11228 13142 11240
rect 13630 11228 13636 11240
rect 13688 11268 13694 11280
rect 14752 11268 14780 11296
rect 13688 11240 14780 11268
rect 13688 11228 13694 11240
rect 14292 11209 14320 11240
rect 14277 11203 14335 11209
rect 13004 11172 13308 11200
rect 11882 11132 11888 11144
rect 11204 11104 11744 11132
rect 11843 11104 11888 11132
rect 11204 11092 11210 11104
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12039 11135 12097 11141
rect 12039 11101 12051 11135
rect 12085 11132 12097 11135
rect 12158 11132 12164 11144
rect 12085 11104 12164 11132
rect 12085 11101 12097 11104
rect 12039 11095 12097 11101
rect 12158 11092 12164 11104
rect 12216 11092 12222 11144
rect 12894 11132 12900 11144
rect 12855 11104 12900 11132
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 12986 11092 12992 11144
rect 13044 11132 13050 11144
rect 13280 11141 13308 11172
rect 14277 11169 14289 11203
rect 14323 11169 14335 11203
rect 14277 11163 14335 11169
rect 14550 11160 14556 11212
rect 14608 11200 14614 11212
rect 14737 11203 14795 11209
rect 14737 11200 14749 11203
rect 14608 11172 14749 11200
rect 14608 11160 14614 11172
rect 14737 11169 14749 11172
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 13265 11135 13323 11141
rect 13044 11104 13089 11132
rect 13044 11092 13050 11104
rect 13265 11101 13277 11135
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 14369 11135 14427 11141
rect 14369 11101 14381 11135
rect 14415 11132 14427 11135
rect 14645 11135 14703 11141
rect 14645 11132 14657 11135
rect 14415 11104 14657 11132
rect 14415 11101 14427 11104
rect 14369 11095 14427 11101
rect 14645 11101 14657 11104
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 7466 11064 7472 11076
rect 6840 11036 7472 11064
rect 7466 11024 7472 11036
rect 7524 11024 7530 11076
rect 7558 11024 7564 11076
rect 7616 11064 7622 11076
rect 7926 11064 7932 11076
rect 7616 11036 7932 11064
rect 7616 11024 7622 11036
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 8772 11036 9076 11064
rect 4522 10956 4528 11008
rect 4580 10996 4586 11008
rect 5445 10999 5503 11005
rect 5445 10996 5457 10999
rect 4580 10968 5457 10996
rect 4580 10956 4586 10968
rect 5445 10965 5457 10968
rect 5491 10996 5503 10999
rect 7098 10996 7104 11008
rect 5491 10968 7104 10996
rect 5491 10965 5503 10968
rect 5445 10959 5503 10965
rect 7098 10956 7104 10968
rect 7156 10996 7162 11008
rect 8772 10996 8800 11036
rect 8938 10996 8944 11008
rect 7156 10968 8800 10996
rect 8899 10968 8944 10996
rect 7156 10956 7162 10968
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 9048 10996 9076 11036
rect 9306 11024 9312 11076
rect 9364 11064 9370 11076
rect 9861 11067 9919 11073
rect 9861 11064 9873 11067
rect 9364 11036 9873 11064
rect 9364 11024 9370 11036
rect 9861 11033 9873 11036
rect 9907 11033 9919 11067
rect 10042 11064 10048 11076
rect 10003 11036 10048 11064
rect 9861 11027 9919 11033
rect 10042 11024 10048 11036
rect 10100 11024 10106 11076
rect 10226 11024 10232 11076
rect 10284 11064 10290 11076
rect 10502 11064 10508 11076
rect 10284 11036 10508 11064
rect 10284 11024 10290 11036
rect 10502 11024 10508 11036
rect 10560 11064 10566 11076
rect 11425 11067 11483 11073
rect 11425 11064 11437 11067
rect 10560 11036 11437 11064
rect 10560 11024 10566 11036
rect 11425 11033 11437 11036
rect 11471 11064 11483 11067
rect 12434 11064 12440 11076
rect 11471 11036 12440 11064
rect 11471 11033 11483 11036
rect 11425 11027 11483 11033
rect 12434 11024 12440 11036
rect 12492 11024 12498 11076
rect 13004 11064 13032 11092
rect 14384 11064 14412 11095
rect 13004 11036 14412 11064
rect 13906 10996 13912 11008
rect 9048 10968 13912 10996
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 1104 10906 15732 10928
rect 1104 10854 5858 10906
rect 5910 10854 5922 10906
rect 5974 10854 5986 10906
rect 6038 10854 6050 10906
rect 6102 10854 10734 10906
rect 10786 10854 10798 10906
rect 10850 10854 10862 10906
rect 10914 10854 10926 10906
rect 10978 10854 15732 10906
rect 1104 10832 15732 10854
rect 2038 10792 2044 10804
rect 1999 10764 2044 10792
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 3602 10792 3608 10804
rect 3563 10764 3608 10792
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 4341 10795 4399 10801
rect 4341 10761 4353 10795
rect 4387 10792 4399 10795
rect 4890 10792 4896 10804
rect 4387 10764 4896 10792
rect 4387 10761 4399 10764
rect 4341 10755 4399 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 6457 10795 6515 10801
rect 6457 10792 6469 10795
rect 5040 10764 6469 10792
rect 5040 10752 5046 10764
rect 6457 10761 6469 10764
rect 6503 10761 6515 10795
rect 6457 10755 6515 10761
rect 6546 10752 6552 10804
rect 6604 10792 6610 10804
rect 6822 10792 6828 10804
rect 6604 10764 6828 10792
rect 6604 10752 6610 10764
rect 6822 10752 6828 10764
rect 6880 10792 6886 10804
rect 7282 10792 7288 10804
rect 6880 10764 7288 10792
rect 6880 10752 6886 10764
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 9122 10752 9128 10804
rect 9180 10792 9186 10804
rect 9217 10795 9275 10801
rect 9217 10792 9229 10795
rect 9180 10764 9229 10792
rect 9180 10752 9186 10764
rect 9217 10761 9229 10764
rect 9263 10761 9275 10795
rect 9217 10755 9275 10761
rect 12066 10752 12072 10804
rect 12124 10792 12130 10804
rect 12124 10764 14596 10792
rect 12124 10752 12130 10764
rect 4157 10727 4215 10733
rect 4157 10724 4169 10727
rect 3528 10696 4169 10724
rect 2222 10656 2228 10668
rect 2183 10628 2228 10656
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2498 10656 2504 10668
rect 2363 10628 2504 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10625 2651 10659
rect 2593 10619 2651 10625
rect 2406 10548 2412 10600
rect 2464 10588 2470 10600
rect 2608 10588 2636 10619
rect 3234 10616 3240 10668
rect 3292 10656 3298 10668
rect 3528 10665 3556 10696
rect 4157 10693 4169 10696
rect 4203 10693 4215 10727
rect 4157 10687 4215 10693
rect 4433 10727 4491 10733
rect 4433 10693 4445 10727
rect 4479 10724 4491 10727
rect 5350 10724 5356 10736
rect 4479 10696 5356 10724
rect 4479 10693 4491 10696
rect 4433 10687 4491 10693
rect 5350 10684 5356 10696
rect 5408 10684 5414 10736
rect 5445 10727 5503 10733
rect 5445 10693 5457 10727
rect 5491 10724 5503 10727
rect 5534 10724 5540 10736
rect 5491 10696 5540 10724
rect 5491 10693 5503 10696
rect 5445 10687 5503 10693
rect 5534 10684 5540 10696
rect 5592 10724 5598 10736
rect 9030 10724 9036 10736
rect 5592 10696 6408 10724
rect 5592 10684 5598 10696
rect 3513 10659 3571 10665
rect 3513 10656 3525 10659
rect 3292 10628 3525 10656
rect 3292 10616 3298 10628
rect 3513 10625 3525 10628
rect 3559 10625 3571 10659
rect 3513 10619 3571 10625
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10625 3755 10659
rect 4522 10656 4528 10668
rect 4483 10628 4528 10656
rect 3697 10619 3755 10625
rect 2464 10560 2636 10588
rect 3712 10588 3740 10619
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 5718 10656 5724 10668
rect 5675 10628 5724 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 6380 10665 6408 10696
rect 6564 10696 9036 10724
rect 6564 10665 6592 10696
rect 9030 10684 9036 10696
rect 9088 10684 9094 10736
rect 9766 10724 9772 10736
rect 9508 10696 9772 10724
rect 6365 10659 6423 10665
rect 6365 10625 6377 10659
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10625 6607 10659
rect 7190 10656 7196 10668
rect 7151 10628 7196 10656
rect 6549 10619 6607 10625
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10656 7619 10659
rect 7834 10656 7840 10668
rect 7607 10628 7840 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 7009 10591 7067 10597
rect 7009 10588 7021 10591
rect 3712 10560 7021 10588
rect 2464 10548 2470 10560
rect 7009 10557 7021 10560
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 4614 10480 4620 10532
rect 4672 10520 4678 10532
rect 4709 10523 4767 10529
rect 4709 10520 4721 10523
rect 4672 10492 4721 10520
rect 4672 10480 4678 10492
rect 4709 10489 4721 10492
rect 4755 10489 4767 10523
rect 4709 10483 4767 10489
rect 5813 10523 5871 10529
rect 5813 10489 5825 10523
rect 5859 10520 5871 10523
rect 6730 10520 6736 10532
rect 5859 10492 6736 10520
rect 5859 10489 5871 10492
rect 5813 10483 5871 10489
rect 6730 10480 6736 10492
rect 6788 10480 6794 10532
rect 7300 10520 7328 10619
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10656 8079 10659
rect 8297 10659 8355 10665
rect 8067 10628 8248 10656
rect 8067 10625 8079 10628
rect 8021 10619 8079 10625
rect 7466 10588 7472 10600
rect 7379 10560 7472 10588
rect 7466 10548 7472 10560
rect 7524 10588 7530 10600
rect 8036 10588 8064 10619
rect 7524 10560 8064 10588
rect 8113 10591 8171 10597
rect 7524 10548 7530 10560
rect 8113 10557 8125 10591
rect 8159 10557 8171 10591
rect 8220 10588 8248 10628
rect 8297 10625 8309 10659
rect 8343 10656 8355 10659
rect 8938 10656 8944 10668
rect 8343 10628 8944 10656
rect 8343 10625 8355 10628
rect 8297 10619 8355 10625
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9508 10665 9536 10696
rect 9766 10684 9772 10696
rect 9824 10684 9830 10736
rect 10410 10684 10416 10736
rect 10468 10724 10474 10736
rect 10505 10727 10563 10733
rect 10505 10724 10517 10727
rect 10468 10696 10517 10724
rect 10468 10684 10474 10696
rect 10505 10693 10517 10696
rect 10551 10693 10563 10727
rect 10505 10687 10563 10693
rect 11974 10684 11980 10736
rect 12032 10724 12038 10736
rect 12032 10696 13032 10724
rect 12032 10684 12038 10696
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 9582 10616 9588 10668
rect 9640 10656 9646 10668
rect 9640 10628 10456 10656
rect 9640 10616 9646 10628
rect 9401 10591 9459 10597
rect 8220 10560 8892 10588
rect 8113 10551 8171 10557
rect 7558 10520 7564 10532
rect 7300 10492 7564 10520
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 7926 10480 7932 10532
rect 7984 10520 7990 10532
rect 8128 10520 8156 10551
rect 8864 10520 8892 10560
rect 9401 10557 9413 10591
rect 9447 10588 9459 10591
rect 9858 10588 9864 10600
rect 9447 10560 9864 10588
rect 9447 10557 9459 10560
rect 9401 10551 9459 10557
rect 9858 10548 9864 10560
rect 9916 10588 9922 10600
rect 10321 10591 10379 10597
rect 10321 10588 10333 10591
rect 9916 10560 10333 10588
rect 9916 10548 9922 10560
rect 10321 10557 10333 10560
rect 10367 10557 10379 10591
rect 10428 10588 10456 10628
rect 10686 10616 10692 10668
rect 10744 10656 10750 10668
rect 11701 10659 11759 10665
rect 10744 10628 10789 10656
rect 10744 10616 10750 10628
rect 11701 10625 11713 10659
rect 11747 10656 11759 10659
rect 12066 10656 12072 10668
rect 11747 10628 12072 10656
rect 11747 10625 11759 10628
rect 11701 10619 11759 10625
rect 12066 10616 12072 10628
rect 12124 10656 12130 10668
rect 12437 10659 12495 10665
rect 12437 10656 12449 10659
rect 12124 10628 12449 10656
rect 12124 10616 12130 10628
rect 12437 10625 12449 10628
rect 12483 10625 12495 10659
rect 12437 10619 12495 10625
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10656 12587 10659
rect 12710 10656 12716 10668
rect 12575 10628 12716 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 13004 10665 13032 10696
rect 13078 10684 13084 10736
rect 13136 10724 13142 10736
rect 14568 10733 14596 10764
rect 13909 10727 13967 10733
rect 13909 10724 13921 10727
rect 13136 10696 13921 10724
rect 13136 10684 13142 10696
rect 13909 10693 13921 10696
rect 13955 10693 13967 10727
rect 13909 10687 13967 10693
rect 14553 10727 14611 10733
rect 14553 10693 14565 10727
rect 14599 10693 14611 10727
rect 14553 10687 14611 10693
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10625 13231 10659
rect 13722 10656 13728 10668
rect 13683 10628 13728 10656
rect 13173 10619 13231 10625
rect 10428 10560 12572 10588
rect 10321 10551 10379 10557
rect 12544 10520 12572 10560
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 13188 10588 13216 10619
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 13924 10656 13952 10687
rect 14642 10656 14648 10668
rect 13924 10628 14648 10656
rect 14642 10616 14648 10628
rect 14700 10616 14706 10668
rect 12676 10560 13216 10588
rect 12676 10548 12682 10560
rect 13906 10548 13912 10600
rect 13964 10588 13970 10600
rect 14369 10591 14427 10597
rect 14369 10588 14381 10591
rect 13964 10560 14381 10588
rect 13964 10548 13970 10560
rect 14369 10557 14381 10560
rect 14415 10557 14427 10591
rect 14369 10551 14427 10557
rect 13078 10520 13084 10532
rect 7984 10492 8800 10520
rect 8864 10492 12434 10520
rect 12544 10492 13084 10520
rect 7984 10480 7990 10492
rect 2501 10455 2559 10461
rect 2501 10421 2513 10455
rect 2547 10452 2559 10455
rect 2682 10452 2688 10464
rect 2547 10424 2688 10452
rect 2547 10421 2559 10424
rect 2501 10415 2559 10421
rect 2682 10412 2688 10424
rect 2740 10412 2746 10464
rect 8110 10452 8116 10464
rect 8071 10424 8116 10452
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 8481 10455 8539 10461
rect 8481 10421 8493 10455
rect 8527 10452 8539 10455
rect 8662 10452 8668 10464
rect 8527 10424 8668 10452
rect 8527 10421 8539 10424
rect 8481 10415 8539 10421
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 8772 10452 8800 10492
rect 10594 10452 10600 10464
rect 8772 10424 10600 10452
rect 10594 10412 10600 10424
rect 10652 10412 10658 10464
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 12406 10452 12434 10492
rect 13078 10480 13084 10492
rect 13136 10480 13142 10532
rect 13173 10523 13231 10529
rect 13173 10489 13185 10523
rect 13219 10520 13231 10523
rect 14734 10520 14740 10532
rect 13219 10492 14740 10520
rect 13219 10489 13231 10492
rect 13173 10483 13231 10489
rect 14734 10480 14740 10492
rect 14792 10480 14798 10532
rect 13722 10452 13728 10464
rect 12406 10424 13728 10452
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 1104 10362 15732 10384
rect 1104 10310 3420 10362
rect 3472 10310 3484 10362
rect 3536 10310 3548 10362
rect 3600 10310 3612 10362
rect 3664 10310 8296 10362
rect 8348 10310 8360 10362
rect 8412 10310 8424 10362
rect 8476 10310 8488 10362
rect 8540 10310 13172 10362
rect 13224 10310 13236 10362
rect 13288 10310 13300 10362
rect 13352 10310 13364 10362
rect 13416 10310 15732 10362
rect 1104 10288 15732 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 3145 10251 3203 10257
rect 3145 10217 3157 10251
rect 3191 10248 3203 10251
rect 3970 10248 3976 10260
rect 3191 10220 3976 10248
rect 3191 10217 3203 10220
rect 3145 10211 3203 10217
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 4065 10251 4123 10257
rect 4065 10217 4077 10251
rect 4111 10248 4123 10251
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 4111 10220 7849 10248
rect 4111 10217 4123 10220
rect 4065 10211 4123 10217
rect 7837 10217 7849 10220
rect 7883 10248 7895 10251
rect 8846 10248 8852 10260
rect 7883 10220 8852 10248
rect 7883 10217 7895 10220
rect 7837 10211 7895 10217
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 10042 10208 10048 10260
rect 10100 10248 10106 10260
rect 10781 10251 10839 10257
rect 10781 10248 10793 10251
rect 10100 10220 10793 10248
rect 10100 10208 10106 10220
rect 10781 10217 10793 10220
rect 10827 10217 10839 10251
rect 10781 10211 10839 10217
rect 11882 10208 11888 10260
rect 11940 10248 11946 10260
rect 11977 10251 12035 10257
rect 11977 10248 11989 10251
rect 11940 10220 11989 10248
rect 11940 10208 11946 10220
rect 11977 10217 11989 10220
rect 12023 10217 12035 10251
rect 11977 10211 12035 10217
rect 12158 10208 12164 10260
rect 12216 10248 12222 10260
rect 12986 10248 12992 10260
rect 12216 10220 12992 10248
rect 12216 10208 12222 10220
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13173 10251 13231 10257
rect 13173 10217 13185 10251
rect 13219 10217 13231 10251
rect 13173 10211 13231 10217
rect 2866 10180 2872 10192
rect 1964 10152 2872 10180
rect 1964 10053 1992 10152
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 4430 10140 4436 10192
rect 4488 10180 4494 10192
rect 8757 10183 8815 10189
rect 8757 10180 8769 10183
rect 4488 10152 8769 10180
rect 4488 10140 4494 10152
rect 8757 10149 8769 10152
rect 8803 10149 8815 10183
rect 8864 10180 8892 10208
rect 11241 10183 11299 10189
rect 11241 10180 11253 10183
rect 8864 10152 11253 10180
rect 8757 10143 8815 10149
rect 11241 10149 11253 10152
rect 11287 10180 11299 10183
rect 12434 10180 12440 10192
rect 11287 10152 11928 10180
rect 12395 10152 12440 10180
rect 11287 10149 11299 10152
rect 11241 10143 11299 10149
rect 11900 10124 11928 10152
rect 12434 10140 12440 10152
rect 12492 10140 12498 10192
rect 13078 10140 13084 10192
rect 13136 10180 13142 10192
rect 13188 10180 13216 10211
rect 13136 10152 13216 10180
rect 13136 10140 13142 10152
rect 14366 10140 14372 10192
rect 14424 10140 14430 10192
rect 2682 10072 2688 10124
rect 2740 10112 2746 10124
rect 4617 10115 4675 10121
rect 4617 10112 4629 10115
rect 2740 10084 4629 10112
rect 2740 10072 2746 10084
rect 4617 10081 4629 10084
rect 4663 10081 4675 10115
rect 9674 10112 9680 10124
rect 4617 10075 4675 10081
rect 5000 10084 9536 10112
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10013 2007 10047
rect 2869 10047 2927 10053
rect 2869 10044 2881 10047
rect 1949 10007 2007 10013
rect 2608 10016 2881 10044
rect 2608 9988 2636 10016
rect 2869 10013 2881 10016
rect 2915 10013 2927 10047
rect 2869 10007 2927 10013
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10013 3019 10047
rect 4154 10044 4160 10056
rect 4115 10016 4160 10044
rect 2961 10007 3019 10013
rect 2222 9936 2228 9988
rect 2280 9976 2286 9988
rect 2501 9979 2559 9985
rect 2501 9976 2513 9979
rect 2280 9948 2513 9976
rect 2280 9936 2286 9948
rect 2501 9945 2513 9948
rect 2547 9945 2559 9979
rect 2501 9939 2559 9945
rect 2516 9908 2544 9939
rect 2590 9936 2596 9988
rect 2648 9976 2654 9988
rect 2976 9976 3004 10007
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 4890 10053 4896 10056
rect 4861 10047 4896 10053
rect 4861 10013 4873 10047
rect 4861 10007 4896 10013
rect 4890 10004 4896 10007
rect 4948 10004 4954 10056
rect 5000 10053 5028 10084
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 5537 10047 5595 10053
rect 5537 10044 5549 10047
rect 5491 10016 5549 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5537 10013 5549 10016
rect 5583 10044 5595 10047
rect 5626 10044 5632 10056
rect 5583 10016 5632 10044
rect 5583 10013 5595 10016
rect 5537 10007 5595 10013
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10044 6699 10047
rect 7650 10044 7656 10056
rect 6687 10016 7656 10044
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 7742 10004 7748 10056
rect 7800 10044 7806 10056
rect 7837 10047 7895 10053
rect 7837 10044 7849 10047
rect 7800 10016 7849 10044
rect 7800 10004 7806 10016
rect 7837 10013 7849 10016
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 8110 10044 8116 10056
rect 7984 10016 8029 10044
rect 8071 10016 8116 10044
rect 7984 10004 7990 10016
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 8757 10047 8815 10053
rect 8757 10013 8769 10047
rect 8803 10044 8815 10047
rect 9125 10047 9183 10053
rect 9125 10044 9137 10047
rect 8803 10016 9137 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 9125 10013 9137 10016
rect 9171 10013 9183 10047
rect 9306 10044 9312 10056
rect 9267 10016 9312 10044
rect 9125 10007 9183 10013
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 6273 9979 6331 9985
rect 6273 9976 6285 9979
rect 2648 9948 2693 9976
rect 2746 9948 6285 9976
rect 2648 9936 2654 9948
rect 2746 9908 2774 9948
rect 6273 9945 6285 9948
rect 6319 9945 6331 9979
rect 6273 9939 6331 9945
rect 6457 9979 6515 9985
rect 6457 9945 6469 9979
rect 6503 9976 6515 9979
rect 6546 9976 6552 9988
rect 6503 9948 6552 9976
rect 6503 9945 6515 9948
rect 6457 9939 6515 9945
rect 6546 9936 6552 9948
rect 6604 9936 6610 9988
rect 7006 9976 7012 9988
rect 6840 9948 7012 9976
rect 2516 9880 2774 9908
rect 4614 9868 4620 9920
rect 4672 9908 4678 9920
rect 5445 9911 5503 9917
rect 5445 9908 5457 9911
rect 4672 9880 5457 9908
rect 4672 9868 4678 9880
rect 5445 9877 5457 9880
rect 5491 9877 5503 9911
rect 5445 9871 5503 9877
rect 5629 9911 5687 9917
rect 5629 9877 5641 9911
rect 5675 9908 5687 9911
rect 6840 9908 6868 9948
rect 7006 9936 7012 9948
rect 7064 9936 7070 9988
rect 7282 9936 7288 9988
rect 7340 9976 7346 9988
rect 9030 9976 9036 9988
rect 7340 9948 9036 9976
rect 7340 9936 7346 9948
rect 9030 9936 9036 9948
rect 9088 9936 9094 9988
rect 9508 9976 9536 10084
rect 9600 10084 9680 10112
rect 9600 10053 9628 10084
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 10980 10084 11744 10112
rect 9585 10047 9643 10053
rect 9585 10013 9597 10047
rect 9631 10013 9643 10047
rect 9585 10007 9643 10013
rect 9769 10047 9827 10053
rect 9769 10013 9781 10047
rect 9815 10044 9827 10047
rect 9858 10044 9864 10056
rect 9815 10016 9864 10044
rect 9815 10013 9827 10016
rect 9769 10007 9827 10013
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 10980 10053 11008 10084
rect 11716 10056 11744 10084
rect 11882 10072 11888 10124
rect 11940 10072 11946 10124
rect 14093 10115 14151 10121
rect 14093 10081 14105 10115
rect 14139 10112 14151 10115
rect 14384 10112 14412 10140
rect 14139 10084 14412 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 10965 10047 11023 10053
rect 10965 10013 10977 10047
rect 11011 10013 11023 10047
rect 10965 10007 11023 10013
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11333 10047 11391 10053
rect 11112 10016 11157 10044
rect 11112 10004 11118 10016
rect 11333 10013 11345 10047
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11348 9976 11376 10007
rect 11698 10004 11704 10056
rect 11756 10044 11762 10056
rect 12158 10044 12164 10056
rect 11756 10016 12164 10044
rect 11756 10004 11762 10016
rect 12158 10004 12164 10016
rect 12216 10004 12222 10056
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 11790 9976 11796 9988
rect 9508 9948 10456 9976
rect 11348 9948 11796 9976
rect 5675 9880 6868 9908
rect 5675 9877 5687 9880
rect 5629 9871 5687 9877
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7653 9911 7711 9917
rect 7653 9908 7665 9911
rect 6972 9880 7665 9908
rect 6972 9868 6978 9880
rect 7653 9877 7665 9880
rect 7699 9877 7711 9911
rect 7653 9871 7711 9877
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 10226 9908 10232 9920
rect 7800 9880 10232 9908
rect 7800 9868 7806 9880
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 10428 9908 10456 9948
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 11882 9936 11888 9988
rect 11940 9976 11946 9988
rect 12268 9976 12296 10007
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 12529 10047 12587 10053
rect 12529 10044 12541 10047
rect 12492 10016 12541 10044
rect 12492 10004 12498 10016
rect 12529 10013 12541 10016
rect 12575 10013 12587 10047
rect 12529 10007 12587 10013
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 11940 9948 12296 9976
rect 11940 9936 11946 9948
rect 11238 9908 11244 9920
rect 10428 9880 11244 9908
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 12268 9908 12296 9948
rect 12989 9979 13047 9985
rect 12989 9945 13001 9979
rect 13035 9945 13047 9979
rect 13188 9976 13216 10007
rect 13262 10004 13268 10056
rect 13320 10044 13326 10056
rect 13320 10016 13365 10044
rect 13320 10004 13326 10016
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 14369 10047 14427 10053
rect 14369 10044 14381 10047
rect 13780 10016 14381 10044
rect 13780 10004 13786 10016
rect 14369 10013 14381 10016
rect 14415 10013 14427 10047
rect 14369 10007 14427 10013
rect 13354 9976 13360 9988
rect 13188 9948 13360 9976
rect 12989 9939 13047 9945
rect 13004 9908 13032 9939
rect 13354 9936 13360 9948
rect 13412 9936 13418 9988
rect 12268 9880 13032 9908
rect 13078 9868 13084 9920
rect 13136 9908 13142 9920
rect 13449 9911 13507 9917
rect 13449 9908 13461 9911
rect 13136 9880 13461 9908
rect 13136 9868 13142 9880
rect 13449 9877 13461 9880
rect 13495 9877 13507 9911
rect 13449 9871 13507 9877
rect 1104 9818 15732 9840
rect 1104 9766 5858 9818
rect 5910 9766 5922 9818
rect 5974 9766 5986 9818
rect 6038 9766 6050 9818
rect 6102 9766 10734 9818
rect 10786 9766 10798 9818
rect 10850 9766 10862 9818
rect 10914 9766 10926 9818
rect 10978 9766 15732 9818
rect 1104 9744 15732 9766
rect 2041 9707 2099 9713
rect 2041 9673 2053 9707
rect 2087 9704 2099 9707
rect 2590 9704 2596 9716
rect 2087 9676 2596 9704
rect 2087 9673 2099 9676
rect 2041 9667 2099 9673
rect 2590 9664 2596 9676
rect 2648 9664 2654 9716
rect 4154 9664 4160 9716
rect 4212 9704 4218 9716
rect 6362 9704 6368 9716
rect 4212 9676 6368 9704
rect 4212 9664 4218 9676
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 6748 9676 8156 9704
rect 2682 9636 2688 9648
rect 2608 9608 2688 9636
rect 2608 9577 2636 9608
rect 2682 9596 2688 9608
rect 2740 9596 2746 9648
rect 3988 9608 4476 9636
rect 3988 9577 4016 9608
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9568 2375 9571
rect 2593 9571 2651 9577
rect 2593 9568 2605 9571
rect 2363 9540 2605 9568
rect 2363 9537 2375 9540
rect 2317 9531 2375 9537
rect 2593 9537 2605 9540
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 3973 9571 4031 9577
rect 3973 9537 3985 9571
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9568 4123 9571
rect 4111 9540 4384 9568
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9500 2283 9503
rect 2406 9500 2412 9512
rect 2271 9472 2412 9500
rect 2271 9469 2283 9472
rect 2225 9463 2283 9469
rect 2406 9460 2412 9472
rect 2464 9500 2470 9512
rect 4356 9509 4384 9540
rect 4448 9512 4476 9608
rect 4982 9596 4988 9648
rect 5040 9636 5046 9648
rect 6748 9636 6776 9676
rect 8128 9674 8156 9676
rect 8128 9646 8248 9674
rect 9306 9664 9312 9716
rect 9364 9704 9370 9716
rect 9493 9707 9551 9713
rect 9493 9704 9505 9707
rect 9364 9676 9505 9704
rect 9364 9664 9370 9676
rect 9493 9673 9505 9676
rect 9539 9673 9551 9707
rect 9493 9667 9551 9673
rect 9582 9664 9588 9716
rect 9640 9704 9646 9716
rect 9861 9707 9919 9713
rect 9861 9704 9873 9707
rect 9640 9676 9873 9704
rect 9640 9664 9646 9676
rect 9861 9673 9873 9676
rect 9907 9673 9919 9707
rect 9861 9667 9919 9673
rect 10410 9664 10416 9716
rect 10468 9704 10474 9716
rect 10597 9707 10655 9713
rect 10597 9704 10609 9707
rect 10468 9676 10609 9704
rect 10468 9664 10474 9676
rect 10597 9673 10609 9676
rect 10643 9673 10655 9707
rect 10597 9667 10655 9673
rect 11146 9664 11152 9716
rect 11204 9704 11210 9716
rect 11609 9707 11667 9713
rect 11609 9704 11621 9707
rect 11204 9676 11621 9704
rect 11204 9664 11210 9676
rect 11609 9673 11621 9676
rect 11655 9673 11667 9707
rect 11609 9667 11667 9673
rect 11790 9664 11796 9716
rect 11848 9704 11854 9716
rect 12434 9704 12440 9716
rect 11848 9676 12440 9704
rect 11848 9664 11854 9676
rect 12434 9664 12440 9676
rect 12492 9704 12498 9716
rect 12802 9704 12808 9716
rect 12492 9676 12808 9704
rect 12492 9664 12498 9676
rect 12802 9664 12808 9676
rect 12860 9704 12866 9716
rect 13262 9704 13268 9716
rect 12860 9676 13268 9704
rect 12860 9664 12866 9676
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 5040 9608 5580 9636
rect 5040 9596 5046 9608
rect 5092 9577 5120 9608
rect 5552 9577 5580 9608
rect 6656 9608 6776 9636
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9537 5227 9571
rect 5169 9531 5227 9537
rect 5537 9571 5595 9577
rect 5537 9537 5549 9571
rect 5583 9568 5595 9571
rect 5626 9568 5632 9580
rect 5583 9540 5632 9568
rect 5583 9537 5595 9540
rect 5537 9531 5595 9537
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2464 9472 2697 9500
rect 2464 9460 2470 9472
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9469 4399 9503
rect 4341 9463 4399 9469
rect 2700 9364 2728 9463
rect 2958 9392 2964 9444
rect 3016 9432 3022 9444
rect 3789 9435 3847 9441
rect 3789 9432 3801 9435
rect 3016 9404 3801 9432
rect 3016 9392 3022 9404
rect 3789 9401 3801 9404
rect 3835 9401 3847 9435
rect 4356 9432 4384 9463
rect 4430 9460 4436 9512
rect 4488 9500 4494 9512
rect 5184 9500 5212 9531
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 5718 9528 5724 9580
rect 5776 9568 5782 9580
rect 6656 9568 6684 9608
rect 7006 9577 7012 9580
rect 5776 9540 6684 9568
rect 6826 9571 6884 9577
rect 5776 9528 5782 9540
rect 6826 9537 6838 9571
rect 6872 9537 6884 9571
rect 6826 9531 6884 9537
rect 6977 9571 7012 9577
rect 6977 9537 6989 9571
rect 6977 9531 7012 9537
rect 5442 9500 5448 9512
rect 4488 9472 4533 9500
rect 5184 9472 5448 9500
rect 4488 9460 4494 9472
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 6840 9500 6868 9531
rect 7006 9528 7012 9531
rect 7064 9528 7070 9580
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9568 7251 9571
rect 7650 9568 7656 9580
rect 7239 9540 7656 9568
rect 7239 9537 7251 9540
rect 7193 9531 7251 9537
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 7926 9568 7932 9580
rect 7791 9540 7932 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 8220 9568 8248 9646
rect 9677 9639 9735 9645
rect 9677 9605 9689 9639
rect 9723 9605 9735 9639
rect 9677 9599 9735 9605
rect 8220 9540 9628 9568
rect 7282 9500 7288 9512
rect 6840 9472 7288 9500
rect 7282 9460 7288 9472
rect 7340 9500 7346 9512
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7340 9472 8033 9500
rect 7340 9460 7346 9472
rect 8021 9469 8033 9472
rect 8067 9469 8079 9503
rect 8021 9463 8079 9469
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9490 9500 9496 9512
rect 9180 9472 9496 9500
rect 9180 9460 9186 9472
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 4706 9432 4712 9444
rect 4356 9404 4712 9432
rect 3789 9395 3847 9401
rect 4706 9392 4712 9404
rect 4764 9432 4770 9444
rect 4893 9435 4951 9441
rect 4893 9432 4905 9435
rect 4764 9404 4905 9432
rect 4764 9392 4770 9404
rect 4893 9401 4905 9404
rect 4939 9401 4951 9435
rect 9306 9432 9312 9444
rect 4893 9395 4951 9401
rect 6288 9404 9312 9432
rect 6288 9364 6316 9404
rect 9306 9392 9312 9404
rect 9364 9392 9370 9444
rect 2700 9336 6316 9364
rect 6362 9324 6368 9376
rect 6420 9364 6426 9376
rect 6641 9367 6699 9373
rect 6641 9364 6653 9367
rect 6420 9336 6653 9364
rect 6420 9324 6426 9336
rect 6641 9333 6653 9336
rect 6687 9333 6699 9367
rect 6641 9327 6699 9333
rect 7101 9367 7159 9373
rect 7101 9333 7113 9367
rect 7147 9364 7159 9367
rect 7926 9364 7932 9376
rect 7147 9336 7932 9364
rect 7147 9333 7159 9336
rect 7101 9327 7159 9333
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 9600 9364 9628 9540
rect 9692 9512 9720 9599
rect 11882 9596 11888 9648
rect 11940 9636 11946 9648
rect 12069 9639 12127 9645
rect 12069 9636 12081 9639
rect 11940 9608 12081 9636
rect 11940 9596 11946 9608
rect 12069 9605 12081 9608
rect 12115 9605 12127 9639
rect 12069 9599 12127 9605
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9537 9827 9571
rect 9769 9534 9827 9537
rect 9769 9531 9904 9534
rect 9674 9460 9680 9512
rect 9732 9460 9738 9512
rect 9788 9506 9904 9531
rect 10318 9528 10324 9580
rect 10376 9568 10382 9580
rect 10505 9571 10563 9577
rect 10505 9568 10517 9571
rect 10376 9540 10517 9568
rect 10376 9528 10382 9540
rect 10505 9537 10517 9540
rect 10551 9537 10563 9571
rect 11790 9568 11796 9580
rect 11751 9540 11796 9568
rect 10505 9531 10563 9537
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 13265 9571 13323 9577
rect 13265 9568 13277 9571
rect 12860 9540 13277 9568
rect 12860 9528 12866 9540
rect 13265 9537 13277 9540
rect 13311 9537 13323 9571
rect 13265 9531 13323 9537
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 14645 9571 14703 9577
rect 14645 9568 14657 9571
rect 13780 9540 14657 9568
rect 13780 9528 13786 9540
rect 14645 9537 14657 9540
rect 14691 9537 14703 9571
rect 14645 9531 14703 9537
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9568 14795 9571
rect 15102 9568 15108 9580
rect 14783 9540 15108 9568
rect 14783 9537 14795 9540
rect 14737 9531 14795 9537
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 9876 9500 9904 9506
rect 10594 9500 10600 9512
rect 9876 9472 10600 9500
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 11698 9460 11704 9512
rect 11756 9500 11762 9512
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 11756 9472 11897 9500
rect 11756 9460 11762 9472
rect 11885 9469 11897 9472
rect 11931 9469 11943 9503
rect 11885 9463 11943 9469
rect 12342 9460 12348 9512
rect 12400 9500 12406 9512
rect 12894 9500 12900 9512
rect 12400 9472 12900 9500
rect 12400 9460 12406 9472
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 14274 9460 14280 9512
rect 14332 9500 14338 9512
rect 14369 9503 14427 9509
rect 14369 9500 14381 9503
rect 14332 9472 14381 9500
rect 14332 9460 14338 9472
rect 14369 9469 14381 9472
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 14458 9460 14464 9512
rect 14516 9500 14522 9512
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 14516 9472 14565 9500
rect 14516 9460 14522 9472
rect 14553 9469 14565 9472
rect 14599 9469 14611 9503
rect 14553 9463 14611 9469
rect 14826 9460 14832 9512
rect 14884 9500 14890 9512
rect 14884 9472 14929 9500
rect 14884 9460 14890 9472
rect 10045 9435 10103 9441
rect 10045 9401 10057 9435
rect 10091 9432 10103 9435
rect 13814 9432 13820 9444
rect 10091 9404 13820 9432
rect 10091 9401 10103 9404
rect 10045 9395 10103 9401
rect 13814 9392 13820 9404
rect 13872 9392 13878 9444
rect 11054 9364 11060 9376
rect 9600 9336 11060 9364
rect 11054 9324 11060 9336
rect 11112 9364 11118 9376
rect 11793 9367 11851 9373
rect 11793 9364 11805 9367
rect 11112 9336 11805 9364
rect 11112 9324 11118 9336
rect 11793 9333 11805 9336
rect 11839 9333 11851 9367
rect 11793 9327 11851 9333
rect 12250 9324 12256 9376
rect 12308 9364 12314 9376
rect 12986 9364 12992 9376
rect 12308 9336 12992 9364
rect 12308 9324 12314 9336
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 1104 9274 15732 9296
rect 1104 9222 3420 9274
rect 3472 9222 3484 9274
rect 3536 9222 3548 9274
rect 3600 9222 3612 9274
rect 3664 9222 8296 9274
rect 8348 9222 8360 9274
rect 8412 9222 8424 9274
rect 8476 9222 8488 9274
rect 8540 9222 13172 9274
rect 13224 9222 13236 9274
rect 13288 9222 13300 9274
rect 13352 9222 13364 9274
rect 13416 9222 15732 9274
rect 1104 9200 15732 9222
rect 2314 9160 2320 9172
rect 2275 9132 2320 9160
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 4893 9163 4951 9169
rect 4893 9129 4905 9163
rect 4939 9160 4951 9163
rect 5442 9160 5448 9172
rect 4939 9132 5448 9160
rect 4939 9129 4951 9132
rect 4893 9123 4951 9129
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 5813 9163 5871 9169
rect 5813 9129 5825 9163
rect 5859 9160 5871 9163
rect 5997 9163 6055 9169
rect 5997 9160 6009 9163
rect 5859 9132 6009 9160
rect 5859 9129 5871 9132
rect 5813 9123 5871 9129
rect 5997 9129 6009 9132
rect 6043 9129 6055 9163
rect 6362 9160 6368 9172
rect 6323 9132 6368 9160
rect 5997 9123 6055 9129
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 7006 9120 7012 9172
rect 7064 9160 7070 9172
rect 7837 9163 7895 9169
rect 7837 9160 7849 9163
rect 7064 9132 7849 9160
rect 7064 9120 7070 9132
rect 7837 9129 7849 9132
rect 7883 9160 7895 9163
rect 8110 9160 8116 9172
rect 7883 9132 8116 9160
rect 7883 9129 7895 9132
rect 7837 9123 7895 9129
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 8754 9120 8760 9172
rect 8812 9160 8818 9172
rect 9030 9160 9036 9172
rect 8812 9132 9036 9160
rect 8812 9120 8818 9132
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 9306 9160 9312 9172
rect 9267 9132 9312 9160
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 10873 9163 10931 9169
rect 10873 9129 10885 9163
rect 10919 9160 10931 9163
rect 11422 9160 11428 9172
rect 10919 9132 11428 9160
rect 10919 9129 10931 9132
rect 10873 9123 10931 9129
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 12802 9160 12808 9172
rect 11532 9132 11744 9160
rect 12763 9132 12808 9160
rect 3237 9095 3295 9101
rect 3237 9061 3249 9095
rect 3283 9092 3295 9095
rect 11054 9092 11060 9104
rect 3283 9064 11060 9092
rect 3283 9061 3295 9064
rect 3237 9055 3295 9061
rect 11054 9052 11060 9064
rect 11112 9052 11118 9104
rect 11532 9092 11560 9132
rect 11164 9064 11560 9092
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 9024 1731 9027
rect 1719 8996 2176 9024
rect 1719 8993 1731 8996
rect 1673 8987 1731 8993
rect 2148 8968 2176 8996
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 7374 9024 7380 9036
rect 4028 8996 7380 9024
rect 4028 8984 4034 8996
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 7466 8984 7472 9036
rect 7524 9024 7530 9036
rect 11164 9024 11192 9064
rect 7524 8996 7696 9024
rect 7524 8984 7530 8996
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 1872 8928 2053 8956
rect 1872 8900 1900 8928
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 3053 8959 3111 8965
rect 2188 8928 2233 8956
rect 2188 8916 2194 8928
rect 3053 8925 3065 8959
rect 3099 8925 3111 8959
rect 3786 8956 3792 8968
rect 3747 8928 3792 8956
rect 3053 8919 3111 8925
rect 1765 8891 1823 8897
rect 1765 8857 1777 8891
rect 1811 8888 1823 8891
rect 1854 8888 1860 8900
rect 1811 8860 1860 8888
rect 1811 8857 1823 8860
rect 1765 8851 1823 8857
rect 1854 8848 1860 8860
rect 1912 8848 1918 8900
rect 3068 8888 3096 8919
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 4430 8916 4436 8968
rect 4488 8956 4494 8968
rect 4617 8959 4675 8965
rect 4617 8956 4629 8959
rect 4488 8928 4629 8956
rect 4488 8916 4494 8928
rect 4617 8925 4629 8928
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 4632 8888 4660 8919
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 4982 8956 4988 8968
rect 4764 8928 4809 8956
rect 4943 8928 4988 8956
rect 4764 8916 4770 8928
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8956 6515 8959
rect 6914 8956 6920 8968
rect 6503 8928 6920 8956
rect 6503 8925 6515 8928
rect 6457 8919 6515 8925
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 7282 8956 7288 8968
rect 7116 8928 7288 8956
rect 5813 8891 5871 8897
rect 5813 8888 5825 8891
rect 3068 8860 4568 8888
rect 4632 8860 5825 8888
rect 3970 8820 3976 8832
rect 3931 8792 3976 8820
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 4433 8823 4491 8829
rect 4433 8820 4445 8823
rect 4120 8792 4445 8820
rect 4120 8780 4126 8792
rect 4433 8789 4445 8792
rect 4479 8789 4491 8823
rect 4540 8820 4568 8860
rect 5813 8857 5825 8860
rect 5859 8857 5871 8891
rect 5813 8851 5871 8857
rect 6546 8848 6552 8900
rect 6604 8888 6610 8900
rect 7116 8888 7144 8928
rect 7282 8916 7288 8928
rect 7340 8956 7346 8968
rect 7668 8965 7696 8996
rect 7760 8996 11192 9024
rect 11716 9024 11744 9132
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 14458 9160 14464 9172
rect 14419 9132 14464 9160
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 12434 9092 12440 9104
rect 12406 9052 12440 9092
rect 12492 9052 12498 9104
rect 12406 9024 12434 9052
rect 11716 8996 12434 9024
rect 13004 8996 14136 9024
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 7340 8928 7573 8956
rect 7340 8916 7346 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 7760 8888 7788 8996
rect 7926 8956 7932 8968
rect 7887 8928 7932 8956
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 9769 8959 9827 8965
rect 9769 8956 9781 8959
rect 9048 8928 9781 8956
rect 6604 8860 7144 8888
rect 7208 8860 7788 8888
rect 7944 8888 7972 8916
rect 8938 8888 8944 8900
rect 7944 8860 8944 8888
rect 6604 8848 6610 8860
rect 7208 8820 7236 8860
rect 8938 8848 8944 8860
rect 8996 8848 9002 8900
rect 7374 8820 7380 8832
rect 4540 8792 7236 8820
rect 7335 8792 7380 8820
rect 4433 8783 4491 8789
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 7466 8780 7472 8832
rect 7524 8820 7530 8832
rect 9048 8820 9076 8928
rect 9769 8925 9781 8928
rect 9815 8956 9827 8959
rect 9858 8956 9864 8968
rect 9815 8928 9864 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 9858 8916 9864 8928
rect 9916 8916 9922 8968
rect 9953 8959 10011 8965
rect 9953 8925 9965 8959
rect 9999 8956 10011 8959
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 9999 8928 10885 8956
rect 9999 8925 10011 8928
rect 9953 8919 10011 8925
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8956 11207 8959
rect 11422 8956 11428 8968
rect 11195 8928 11428 8956
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 9125 8891 9183 8897
rect 9125 8857 9137 8891
rect 9171 8888 9183 8891
rect 9968 8888 9996 8919
rect 11422 8916 11428 8928
rect 11480 8916 11486 8968
rect 11606 8956 11612 8968
rect 11567 8928 11612 8956
rect 11606 8916 11612 8928
rect 11664 8950 11670 8968
rect 13004 8956 13032 8996
rect 11716 8950 13032 8956
rect 11664 8928 13032 8950
rect 13081 8959 13139 8965
rect 11664 8922 11744 8928
rect 13081 8925 13093 8959
rect 13127 8956 13139 8959
rect 13814 8956 13820 8968
rect 13127 8928 13820 8956
rect 13127 8925 13139 8928
rect 11664 8916 11670 8922
rect 13081 8919 13139 8925
rect 13814 8916 13820 8928
rect 13872 8916 13878 8968
rect 14108 8965 14136 8996
rect 14093 8959 14151 8965
rect 14093 8925 14105 8959
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8956 14335 8959
rect 14366 8956 14372 8968
rect 14323 8928 14372 8956
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 9171 8860 9996 8888
rect 9171 8857 9183 8860
rect 9125 8851 9183 8857
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 11793 8891 11851 8897
rect 11793 8888 11805 8891
rect 10468 8860 11805 8888
rect 10468 8848 10474 8860
rect 11793 8857 11805 8860
rect 11839 8857 11851 8891
rect 15010 8888 15016 8900
rect 11793 8851 11851 8857
rect 11900 8860 15016 8888
rect 7524 8792 9076 8820
rect 7524 8780 7530 8792
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 9861 8823 9919 8829
rect 9861 8820 9873 8823
rect 9640 8792 9873 8820
rect 9640 8780 9646 8792
rect 9861 8789 9873 8792
rect 9907 8789 9919 8823
rect 9861 8783 9919 8789
rect 11057 8823 11115 8829
rect 11057 8789 11069 8823
rect 11103 8820 11115 8823
rect 11900 8820 11928 8860
rect 15010 8848 15016 8860
rect 15068 8848 15074 8900
rect 11103 8792 11928 8820
rect 11103 8789 11115 8792
rect 11057 8783 11115 8789
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 12032 8792 12077 8820
rect 12032 8780 12038 8792
rect 1104 8730 15732 8752
rect 1104 8678 5858 8730
rect 5910 8678 5922 8730
rect 5974 8678 5986 8730
rect 6038 8678 6050 8730
rect 6102 8678 10734 8730
rect 10786 8678 10798 8730
rect 10850 8678 10862 8730
rect 10914 8678 10926 8730
rect 10978 8678 15732 8730
rect 1104 8656 15732 8678
rect 5442 8576 5448 8628
rect 5500 8616 5506 8628
rect 9309 8619 9367 8625
rect 9309 8616 9321 8619
rect 5500 8588 9321 8616
rect 5500 8576 5506 8588
rect 9309 8585 9321 8588
rect 9355 8585 9367 8619
rect 10502 8616 10508 8628
rect 9309 8579 9367 8585
rect 9413 8588 10508 8616
rect 3142 8548 3148 8560
rect 1964 8520 2452 8548
rect 1964 8489 1992 8520
rect 2424 8489 2452 8520
rect 2746 8520 3148 8548
rect 2746 8492 2774 8520
rect 3142 8508 3148 8520
rect 3200 8508 3206 8560
rect 4062 8548 4068 8560
rect 3804 8520 4068 8548
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 2409 8483 2467 8489
rect 2087 8452 2360 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2332 8424 2360 8452
rect 2409 8449 2421 8483
rect 2455 8480 2467 8483
rect 2746 8480 2780 8492
rect 2455 8452 2780 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 3804 8489 3832 8520
rect 4062 8508 4068 8520
rect 4120 8548 4126 8560
rect 4249 8551 4307 8557
rect 4249 8548 4261 8551
rect 4120 8520 4261 8548
rect 4120 8508 4126 8520
rect 4249 8517 4261 8520
rect 4295 8517 4307 8551
rect 5813 8551 5871 8557
rect 5813 8548 5825 8551
rect 4249 8511 4307 8517
rect 5368 8520 5825 8548
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3789 8483 3847 8489
rect 3099 8452 3740 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 2314 8412 2320 8424
rect 2275 8384 2320 8412
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 2866 8344 2872 8356
rect 2827 8316 2872 8344
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 3712 8344 3740 8452
rect 3789 8449 3801 8483
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 5368 8489 5396 8520
rect 5813 8517 5825 8520
rect 5859 8548 5871 8551
rect 6914 8548 6920 8560
rect 5859 8520 6920 8548
rect 5859 8517 5871 8520
rect 5813 8511 5871 8517
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 9214 8548 9220 8560
rect 7024 8520 9220 8548
rect 4157 8483 4215 8489
rect 4157 8480 4169 8483
rect 3936 8452 4169 8480
rect 3936 8440 3942 8452
rect 4157 8449 4169 8452
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8449 5503 8483
rect 5445 8443 5503 8449
rect 5460 8412 5488 8443
rect 6362 8440 6368 8492
rect 6420 8480 6426 8492
rect 6457 8483 6515 8489
rect 6457 8480 6469 8483
rect 6420 8452 6469 8480
rect 6420 8440 6426 8452
rect 6457 8449 6469 8452
rect 6503 8449 6515 8483
rect 6457 8443 6515 8449
rect 5718 8412 5724 8424
rect 5460 8384 5724 8412
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 7024 8412 7052 8520
rect 9214 8508 9220 8520
rect 9272 8508 9278 8560
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8480 7619 8483
rect 8662 8480 8668 8492
rect 7607 8452 8668 8480
rect 7607 8449 7619 8452
rect 7561 8443 7619 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 8938 8480 8944 8492
rect 8895 8452 8944 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 9413 8480 9441 8588
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 11517 8619 11575 8625
rect 11517 8616 11529 8619
rect 11296 8588 11529 8616
rect 11296 8576 11302 8588
rect 11517 8585 11529 8588
rect 11563 8585 11575 8619
rect 11517 8579 11575 8585
rect 13722 8576 13728 8628
rect 13780 8576 13786 8628
rect 14458 8576 14464 8628
rect 14516 8576 14522 8628
rect 14553 8619 14611 8625
rect 14553 8585 14565 8619
rect 14599 8616 14611 8619
rect 15194 8616 15200 8628
rect 14599 8588 15200 8616
rect 14599 8585 14611 8588
rect 14553 8579 14611 8585
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 9861 8551 9919 8557
rect 9861 8548 9873 8551
rect 9646 8520 9873 8548
rect 9646 8492 9674 8520
rect 9861 8517 9873 8520
rect 9907 8517 9919 8551
rect 9861 8511 9919 8517
rect 11054 8508 11060 8560
rect 11112 8548 11118 8560
rect 12986 8548 12992 8560
rect 11112 8520 12992 8548
rect 11112 8508 11118 8520
rect 12986 8508 12992 8520
rect 13044 8508 13050 8560
rect 13740 8548 13768 8576
rect 14476 8548 14504 8576
rect 14737 8551 14795 8557
rect 14737 8548 14749 8551
rect 13740 8520 14412 8548
rect 14476 8520 14749 8548
rect 9582 8480 9588 8492
rect 9048 8452 9441 8480
rect 9543 8452 9588 8480
rect 5828 8384 7052 8412
rect 8573 8415 8631 8421
rect 5828 8344 5856 8384
rect 8573 8381 8585 8415
rect 8619 8412 8631 8415
rect 8754 8412 8760 8424
rect 8619 8384 8760 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 8754 8372 8760 8384
rect 8812 8372 8818 8424
rect 9048 8412 9076 8452
rect 9582 8440 9588 8452
rect 9640 8452 9674 8492
rect 10410 8480 10416 8492
rect 10371 8452 10416 8480
rect 9640 8440 9646 8452
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10594 8480 10600 8492
rect 10555 8452 10600 8480
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 11514 8480 11520 8492
rect 11072 8452 11520 8480
rect 11072 8424 11100 8452
rect 11514 8440 11520 8452
rect 11572 8480 11578 8492
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11572 8452 11713 8480
rect 11572 8440 11578 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8480 12127 8483
rect 12894 8480 12900 8492
rect 12115 8452 12900 8480
rect 12115 8449 12127 8452
rect 12069 8443 12127 8449
rect 9490 8412 9496 8424
rect 8864 8384 9076 8412
rect 9403 8384 9496 8412
rect 3712 8316 5856 8344
rect 5902 8304 5908 8356
rect 5960 8344 5966 8356
rect 7101 8347 7159 8353
rect 7101 8344 7113 8347
rect 5960 8316 7113 8344
rect 5960 8304 5966 8316
rect 7101 8313 7113 8316
rect 7147 8313 7159 8347
rect 8864 8344 8892 8384
rect 9490 8372 9496 8384
rect 9548 8412 9554 8424
rect 9953 8415 10011 8421
rect 9953 8412 9965 8415
rect 9548 8384 9965 8412
rect 9548 8372 9554 8384
rect 9953 8381 9965 8384
rect 9999 8412 10011 8415
rect 10505 8415 10563 8421
rect 10505 8412 10517 8415
rect 9999 8384 10517 8412
rect 9999 8381 10011 8384
rect 9953 8375 10011 8381
rect 10505 8381 10517 8384
rect 10551 8381 10563 8415
rect 10505 8375 10563 8381
rect 11054 8372 11060 8424
rect 11112 8372 11118 8424
rect 11606 8372 11612 8424
rect 11664 8412 11670 8424
rect 11809 8412 11837 8443
rect 11664 8384 11837 8412
rect 11664 8372 11670 8384
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 12084 8412 12112 8443
rect 12894 8440 12900 8452
rect 12952 8480 12958 8492
rect 13081 8483 13139 8489
rect 13081 8480 13093 8483
rect 12952 8452 13093 8480
rect 12952 8440 12958 8452
rect 13081 8449 13093 8452
rect 13127 8449 13139 8483
rect 13081 8443 13139 8449
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8480 13323 8483
rect 13538 8480 13544 8492
rect 13311 8452 13544 8480
rect 13311 8449 13323 8452
rect 13265 8443 13323 8449
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 13725 8483 13783 8489
rect 13725 8449 13737 8483
rect 13771 8449 13783 8483
rect 13725 8443 13783 8449
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8480 13875 8483
rect 14274 8480 14280 8492
rect 13863 8452 14280 8480
rect 13863 8449 13875 8452
rect 13817 8443 13875 8449
rect 11940 8384 12112 8412
rect 11940 8372 11946 8384
rect 12802 8372 12808 8424
rect 12860 8412 12866 8424
rect 13446 8412 13452 8424
rect 12860 8384 13452 8412
rect 12860 8372 12866 8384
rect 13446 8372 13452 8384
rect 13504 8412 13510 8424
rect 13740 8412 13768 8443
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 14384 8480 14412 8520
rect 14737 8517 14749 8520
rect 14783 8517 14795 8551
rect 14737 8511 14795 8517
rect 14461 8483 14519 8489
rect 14461 8480 14473 8483
rect 14384 8452 14473 8480
rect 14461 8449 14473 8452
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 13998 8412 14004 8424
rect 13504 8384 13768 8412
rect 13959 8384 14004 8412
rect 13504 8372 13510 8384
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 7101 8307 7159 8313
rect 7208 8316 8892 8344
rect 1765 8279 1823 8285
rect 1765 8245 1777 8279
rect 1811 8276 1823 8279
rect 1854 8276 1860 8288
rect 1811 8248 1860 8276
rect 1811 8245 1823 8248
rect 1765 8239 1823 8245
rect 1854 8236 1860 8248
rect 1912 8236 1918 8288
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 3605 8279 3663 8285
rect 3605 8276 3617 8279
rect 3200 8248 3617 8276
rect 3200 8236 3206 8248
rect 3605 8245 3617 8248
rect 3651 8245 3663 8279
rect 5166 8276 5172 8288
rect 5127 8248 5172 8276
rect 3605 8239 3663 8245
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 6549 8279 6607 8285
rect 6549 8245 6561 8279
rect 6595 8276 6607 8279
rect 7208 8276 7236 8316
rect 9306 8304 9312 8356
rect 9364 8344 9370 8356
rect 9364 8316 9812 8344
rect 9364 8304 9370 8316
rect 7374 8276 7380 8288
rect 6595 8248 7236 8276
rect 7335 8248 7380 8276
rect 6595 8245 6607 8248
rect 6549 8239 6607 8245
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 9784 8276 9812 8316
rect 9858 8304 9864 8356
rect 9916 8344 9922 8356
rect 11977 8347 12035 8353
rect 11977 8344 11989 8347
rect 9916 8316 11989 8344
rect 9916 8304 9922 8316
rect 11977 8313 11989 8316
rect 12023 8313 12035 8347
rect 11977 8307 12035 8313
rect 13909 8347 13967 8353
rect 13909 8313 13921 8347
rect 13955 8344 13967 8347
rect 14550 8344 14556 8356
rect 13955 8316 14556 8344
rect 13955 8313 13967 8316
rect 13909 8307 13967 8313
rect 14550 8304 14556 8316
rect 14608 8304 14614 8356
rect 14737 8347 14795 8353
rect 14737 8313 14749 8347
rect 14783 8344 14795 8347
rect 14826 8344 14832 8356
rect 14783 8316 14832 8344
rect 14783 8313 14795 8316
rect 14737 8307 14795 8313
rect 14826 8304 14832 8316
rect 14884 8304 14890 8356
rect 9950 8276 9956 8288
rect 9784 8248 9956 8276
rect 9950 8236 9956 8248
rect 10008 8236 10014 8288
rect 10686 8236 10692 8288
rect 10744 8276 10750 8288
rect 12710 8276 12716 8288
rect 10744 8248 12716 8276
rect 10744 8236 10750 8248
rect 12710 8236 12716 8248
rect 12768 8236 12774 8288
rect 12894 8276 12900 8288
rect 12855 8248 12900 8276
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 1104 8186 15732 8208
rect 1104 8134 3420 8186
rect 3472 8134 3484 8186
rect 3536 8134 3548 8186
rect 3600 8134 3612 8186
rect 3664 8134 8296 8186
rect 8348 8134 8360 8186
rect 8412 8134 8424 8186
rect 8476 8134 8488 8186
rect 8540 8134 13172 8186
rect 13224 8134 13236 8186
rect 13288 8134 13300 8186
rect 13352 8134 13364 8186
rect 13416 8134 15732 8186
rect 1104 8112 15732 8134
rect 2041 8075 2099 8081
rect 2041 8041 2053 8075
rect 2087 8072 2099 8075
rect 2314 8072 2320 8084
rect 2087 8044 2320 8072
rect 2087 8041 2099 8044
rect 2041 8035 2099 8041
rect 2314 8032 2320 8044
rect 2372 8072 2378 8084
rect 2593 8075 2651 8081
rect 2593 8072 2605 8075
rect 2372 8044 2605 8072
rect 2372 8032 2378 8044
rect 2593 8041 2605 8044
rect 2639 8041 2651 8075
rect 2593 8035 2651 8041
rect 3973 8075 4031 8081
rect 3973 8041 3985 8075
rect 4019 8072 4031 8075
rect 10502 8072 10508 8084
rect 4019 8044 10508 8072
rect 4019 8041 4031 8044
rect 3973 8035 4031 8041
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 10652 8044 10885 8072
rect 10652 8032 10658 8044
rect 10873 8041 10885 8044
rect 10919 8041 10931 8075
rect 12621 8075 12679 8081
rect 12621 8072 12633 8075
rect 10873 8035 10931 8041
rect 12406 8044 12633 8072
rect 3694 8004 3700 8016
rect 2792 7976 3700 8004
rect 2792 7945 2820 7976
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7905 2835 7939
rect 3142 7936 3148 7948
rect 3103 7908 3148 7936
rect 2777 7899 2835 7905
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 3252 7945 3280 7976
rect 3694 7964 3700 7976
rect 3752 8004 3758 8016
rect 4433 8007 4491 8013
rect 4433 8004 4445 8007
rect 3752 7976 4445 8004
rect 3752 7964 3758 7976
rect 4433 7973 4445 7976
rect 4479 7973 4491 8007
rect 4433 7967 4491 7973
rect 4908 7976 5672 8004
rect 3237 7939 3295 7945
rect 3237 7905 3249 7939
rect 3283 7905 3295 7939
rect 4908 7936 4936 7976
rect 3237 7899 3295 7905
rect 3804 7908 4936 7936
rect 4985 7939 5043 7945
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 1578 7732 1584 7744
rect 1539 7704 1584 7732
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 1780 7732 1808 7831
rect 1854 7828 1860 7880
rect 1912 7868 1918 7880
rect 2133 7871 2191 7877
rect 1912 7840 1957 7868
rect 1912 7828 1918 7840
rect 2133 7837 2145 7871
rect 2179 7868 2191 7871
rect 2682 7868 2688 7880
rect 2179 7840 2688 7868
rect 2179 7837 2191 7840
rect 2133 7831 2191 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7868 2927 7871
rect 3160 7868 3188 7896
rect 3804 7877 3832 7908
rect 4985 7905 4997 7939
rect 5031 7936 5043 7939
rect 5166 7936 5172 7948
rect 5031 7908 5172 7936
rect 5031 7905 5043 7908
rect 4985 7899 5043 7905
rect 2915 7840 3188 7868
rect 3789 7871 3847 7877
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 3970 7868 3976 7880
rect 3931 7840 3976 7868
rect 3789 7831 3847 7837
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7868 4767 7871
rect 5000 7868 5028 7899
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 4755 7840 5028 7868
rect 5644 7868 5672 7976
rect 5718 7964 5724 8016
rect 5776 8004 5782 8016
rect 9309 8007 9367 8013
rect 9309 8004 9321 8007
rect 5776 7976 9321 8004
rect 5776 7964 5782 7976
rect 9309 7973 9321 7976
rect 9355 7973 9367 8007
rect 9309 7967 9367 7973
rect 10410 7964 10416 8016
rect 10468 8004 10474 8016
rect 12406 8004 12434 8044
rect 12621 8041 12633 8044
rect 12667 8041 12679 8075
rect 12621 8035 12679 8041
rect 10468 7976 12434 8004
rect 13173 8007 13231 8013
rect 10468 7964 10474 7976
rect 13173 7973 13185 8007
rect 13219 8004 13231 8007
rect 13814 8004 13820 8016
rect 13219 7976 13820 8004
rect 13219 7973 13231 7976
rect 13173 7967 13231 7973
rect 13814 7964 13820 7976
rect 13872 7964 13878 8016
rect 6914 7936 6920 7948
rect 6564 7908 6920 7936
rect 6274 7881 6332 7887
rect 5644 7840 6224 7868
rect 6274 7847 6286 7881
rect 6320 7868 6332 7881
rect 6564 7868 6592 7908
rect 6914 7896 6920 7908
rect 6972 7936 6978 7948
rect 10428 7936 10456 7964
rect 6972 7908 7236 7936
rect 6972 7896 6978 7908
rect 6730 7868 6736 7880
rect 6320 7847 6592 7868
rect 6274 7841 6592 7847
rect 6288 7840 6592 7841
rect 6691 7840 6736 7868
rect 4755 7837 4767 7840
rect 4709 7831 4767 7837
rect 4632 7800 4660 7831
rect 5077 7803 5135 7809
rect 5077 7800 5089 7803
rect 3804 7772 4568 7800
rect 4632 7772 5089 7800
rect 2130 7732 2136 7744
rect 1780 7704 2136 7732
rect 2130 7692 2136 7704
rect 2188 7732 2194 7744
rect 3804 7732 3832 7772
rect 2188 7704 3832 7732
rect 4540 7732 4568 7772
rect 5077 7769 5089 7772
rect 5123 7800 5135 7803
rect 5534 7800 5540 7812
rect 5123 7772 5540 7800
rect 5123 7769 5135 7772
rect 5077 7763 5135 7769
rect 5534 7760 5540 7772
rect 5592 7800 5598 7812
rect 5902 7800 5908 7812
rect 5592 7772 5908 7800
rect 5592 7760 5598 7772
rect 5902 7760 5908 7772
rect 5960 7760 5966 7812
rect 6089 7735 6147 7741
rect 6089 7732 6101 7735
rect 4540 7704 6101 7732
rect 2188 7692 2194 7704
rect 6089 7701 6101 7704
rect 6135 7701 6147 7735
rect 6196 7732 6224 7840
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 7208 7877 7236 7908
rect 9324 7908 10456 7936
rect 11333 7939 11391 7945
rect 7193 7871 7251 7877
rect 7193 7837 7205 7871
rect 7239 7837 7251 7871
rect 7558 7868 7564 7880
rect 7193 7831 7251 7837
rect 7392 7840 7564 7868
rect 6270 7760 6276 7812
rect 6328 7800 6334 7812
rect 6365 7803 6423 7809
rect 6365 7800 6377 7803
rect 6328 7772 6377 7800
rect 6328 7760 6334 7772
rect 6365 7769 6377 7772
rect 6411 7769 6423 7803
rect 6365 7763 6423 7769
rect 6454 7760 6460 7812
rect 6512 7800 6518 7812
rect 6595 7803 6653 7809
rect 6512 7772 6557 7800
rect 6512 7760 6518 7772
rect 6595 7769 6607 7803
rect 6641 7800 6653 7803
rect 6822 7800 6828 7812
rect 6641 7772 6828 7800
rect 6641 7769 6653 7772
rect 6595 7763 6653 7769
rect 6822 7760 6828 7772
rect 6880 7800 6886 7812
rect 7285 7803 7343 7809
rect 7285 7800 7297 7803
rect 6880 7772 7297 7800
rect 6880 7760 6886 7772
rect 7285 7769 7297 7772
rect 7331 7769 7343 7803
rect 7285 7763 7343 7769
rect 7392 7732 7420 7840
rect 7558 7828 7564 7840
rect 7616 7868 7622 7880
rect 9324 7877 9352 7908
rect 11333 7905 11345 7939
rect 11379 7936 11391 7939
rect 11698 7936 11704 7948
rect 11379 7908 11704 7936
rect 11379 7905 11391 7908
rect 11333 7899 11391 7905
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 7616 7840 8401 7868
rect 7616 7828 7622 7840
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7837 9367 7871
rect 9582 7868 9588 7880
rect 9543 7840 9588 7868
rect 9309 7831 9367 7837
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 10410 7868 10416 7880
rect 10371 7840 10416 7868
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 11054 7868 11060 7880
rect 11015 7840 11060 7868
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11425 7871 11483 7877
rect 11204 7840 11249 7868
rect 11204 7828 11210 7840
rect 11425 7837 11437 7871
rect 11471 7868 11483 7871
rect 11882 7868 11888 7880
rect 11471 7840 11888 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 11882 7828 11888 7840
rect 11940 7828 11946 7880
rect 11977 7871 12035 7877
rect 11977 7837 11989 7871
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 9490 7800 9496 7812
rect 9451 7772 9496 7800
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 10042 7760 10048 7812
rect 10100 7800 10106 7812
rect 11606 7800 11612 7812
rect 10100 7772 11612 7800
rect 10100 7760 10106 7772
rect 11606 7760 11612 7772
rect 11664 7800 11670 7812
rect 11992 7800 12020 7831
rect 12710 7828 12716 7880
rect 12768 7868 12774 7880
rect 12897 7871 12955 7877
rect 12897 7868 12909 7871
rect 12768 7840 12909 7868
rect 12768 7828 12774 7840
rect 12897 7837 12909 7840
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 13096 7840 13492 7868
rect 11664 7772 12020 7800
rect 11664 7760 11670 7772
rect 12526 7760 12532 7812
rect 12584 7800 12590 7812
rect 12805 7803 12863 7809
rect 12805 7800 12817 7803
rect 12584 7772 12817 7800
rect 12584 7760 12590 7772
rect 12805 7769 12817 7772
rect 12851 7800 12863 7803
rect 13096 7800 13124 7840
rect 12851 7772 13124 7800
rect 13464 7800 13492 7840
rect 13538 7828 13544 7880
rect 13596 7868 13602 7880
rect 14185 7871 14243 7877
rect 14185 7868 14197 7871
rect 13596 7840 14197 7868
rect 13596 7828 13602 7840
rect 14185 7837 14197 7840
rect 14231 7837 14243 7871
rect 14185 7831 14243 7837
rect 14274 7828 14280 7880
rect 14332 7868 14338 7880
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 14332 7840 14473 7868
rect 14332 7828 14338 7840
rect 14461 7837 14473 7840
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 13722 7800 13728 7812
rect 13464 7772 13728 7800
rect 12851 7769 12863 7772
rect 12805 7763 12863 7769
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 6196 7704 7420 7732
rect 6089 7695 6147 7701
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 8205 7735 8263 7741
rect 8205 7732 8217 7735
rect 7524 7704 8217 7732
rect 7524 7692 7530 7704
rect 8205 7701 8217 7704
rect 8251 7701 8263 7735
rect 8205 7695 8263 7701
rect 10321 7735 10379 7741
rect 10321 7701 10333 7735
rect 10367 7732 10379 7735
rect 11330 7732 11336 7744
rect 10367 7704 11336 7732
rect 10367 7701 10379 7704
rect 10321 7695 10379 7701
rect 11330 7692 11336 7704
rect 11388 7692 11394 7744
rect 11698 7692 11704 7744
rect 11756 7732 11762 7744
rect 12161 7735 12219 7741
rect 12161 7732 12173 7735
rect 11756 7704 12173 7732
rect 11756 7692 11762 7704
rect 12161 7701 12173 7704
rect 12207 7701 12219 7735
rect 12986 7732 12992 7744
rect 12947 7704 12992 7732
rect 12161 7695 12219 7701
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 1104 7642 15732 7664
rect 1104 7590 5858 7642
rect 5910 7590 5922 7642
rect 5974 7590 5986 7642
rect 6038 7590 6050 7642
rect 6102 7590 10734 7642
rect 10786 7590 10798 7642
rect 10850 7590 10862 7642
rect 10914 7590 10926 7642
rect 10978 7590 15732 7642
rect 1104 7568 15732 7590
rect 2961 7531 3019 7537
rect 2961 7497 2973 7531
rect 3007 7528 3019 7531
rect 6914 7528 6920 7540
rect 3007 7500 6776 7528
rect 6875 7500 6920 7528
rect 3007 7497 3019 7500
rect 2961 7491 3019 7497
rect 3142 7420 3148 7472
rect 3200 7460 3206 7472
rect 3200 7432 3832 7460
rect 3200 7420 3206 7432
rect 2866 7392 2872 7404
rect 2827 7364 2872 7392
rect 2866 7352 2872 7364
rect 2924 7352 2930 7404
rect 3694 7392 3700 7404
rect 3655 7364 3700 7392
rect 3694 7352 3700 7364
rect 3752 7352 3758 7404
rect 3804 7401 3832 7432
rect 5166 7420 5172 7472
rect 5224 7460 5230 7472
rect 6748 7460 6776 7500
rect 6914 7488 6920 7500
rect 6972 7488 6978 7540
rect 10042 7528 10048 7540
rect 7024 7500 10048 7528
rect 7024 7460 7052 7500
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 10410 7488 10416 7540
rect 10468 7528 10474 7540
rect 13449 7531 13507 7537
rect 10468 7500 13400 7528
rect 10468 7488 10474 7500
rect 7834 7460 7840 7472
rect 5224 7432 5396 7460
rect 6748 7432 7052 7460
rect 7116 7432 7840 7460
rect 5224 7420 5230 7432
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7361 3847 7395
rect 4062 7392 4068 7404
rect 4023 7364 4068 7392
rect 3789 7355 3847 7361
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 5368 7401 5396 7432
rect 5261 7395 5319 7401
rect 5261 7361 5273 7395
rect 5307 7361 5319 7395
rect 5261 7355 5319 7361
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7392 5687 7395
rect 7006 7392 7012 7404
rect 5675 7364 7012 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 3878 7284 3884 7336
rect 3936 7324 3942 7336
rect 3973 7327 4031 7333
rect 3973 7324 3985 7327
rect 3936 7296 3985 7324
rect 3936 7284 3942 7296
rect 3973 7293 3985 7296
rect 4019 7293 4031 7327
rect 5276 7324 5304 7355
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 7116 7401 7144 7432
rect 7834 7420 7840 7432
rect 7892 7420 7898 7472
rect 11882 7460 11888 7472
rect 9646 7432 11888 7460
rect 7101 7395 7159 7401
rect 7101 7361 7113 7395
rect 7147 7361 7159 7395
rect 7101 7355 7159 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7423 7364 7512 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 5534 7324 5540 7336
rect 5276 7296 5540 7324
rect 3973 7287 4031 7293
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 7282 7324 7288 7336
rect 7195 7296 7288 7324
rect 7282 7284 7288 7296
rect 7340 7324 7346 7336
rect 7484 7324 7512 7364
rect 7558 7352 7564 7404
rect 7616 7392 7622 7404
rect 8205 7395 8263 7401
rect 7616 7364 7661 7392
rect 7616 7352 7622 7364
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 9646 7392 9674 7432
rect 11882 7420 11888 7432
rect 11940 7420 11946 7472
rect 12526 7460 12532 7472
rect 12487 7432 12532 7460
rect 12526 7420 12532 7432
rect 12584 7420 12590 7472
rect 12759 7463 12817 7469
rect 12759 7429 12771 7463
rect 12805 7460 12817 7463
rect 12894 7460 12900 7472
rect 12805 7432 12900 7460
rect 12805 7429 12817 7432
rect 12759 7423 12817 7429
rect 12894 7420 12900 7432
rect 12952 7420 12958 7472
rect 13372 7460 13400 7500
rect 13449 7497 13461 7531
rect 13495 7528 13507 7531
rect 13538 7528 13544 7540
rect 13495 7500 13544 7528
rect 13495 7497 13507 7500
rect 13449 7491 13507 7497
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 13372 7432 14228 7460
rect 14200 7404 14228 7432
rect 9171 7364 9674 7392
rect 9769 7395 9827 7401
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 9769 7361 9781 7395
rect 9815 7392 9827 7395
rect 9858 7392 9864 7404
rect 9815 7364 9864 7392
rect 9815 7361 9827 7364
rect 9769 7355 9827 7361
rect 8220 7324 8248 7355
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 10226 7352 10232 7404
rect 10284 7392 10290 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 10284 7364 10333 7392
rect 10284 7352 10290 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 11609 7395 11667 7401
rect 11609 7392 11621 7395
rect 11204 7364 11621 7392
rect 11204 7352 11210 7364
rect 11609 7361 11621 7364
rect 11655 7392 11667 7395
rect 11790 7392 11796 7404
rect 11655 7364 11796 7392
rect 11655 7361 11667 7364
rect 11609 7355 11667 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 12434 7392 12440 7404
rect 12395 7364 12440 7392
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 12621 7395 12679 7401
rect 12621 7361 12633 7395
rect 12667 7392 12679 7395
rect 12667 7364 13032 7392
rect 12667 7361 12679 7364
rect 12621 7355 12679 7361
rect 10962 7324 10968 7336
rect 7340 7296 7420 7324
rect 7484 7296 10968 7324
rect 7340 7284 7346 7296
rect 7193 7259 7251 7265
rect 7193 7225 7205 7259
rect 7239 7225 7251 7259
rect 7392 7256 7420 7296
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11974 7284 11980 7336
rect 12032 7324 12038 7336
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 12032 7296 12909 7324
rect 12032 7284 12038 7296
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 13004 7324 13032 7364
rect 13078 7352 13084 7404
rect 13136 7392 13142 7404
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 13136 7364 13369 7392
rect 13136 7352 13142 7364
rect 13357 7361 13369 7364
rect 13403 7361 13415 7395
rect 14182 7392 14188 7404
rect 14095 7364 14188 7392
rect 13357 7355 13415 7361
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 14458 7392 14464 7404
rect 14419 7364 14464 7392
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 13814 7324 13820 7336
rect 13004 7296 13820 7324
rect 12897 7287 12955 7293
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 13964 7296 14289 7324
rect 13964 7284 13970 7296
rect 14277 7293 14289 7296
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 14366 7284 14372 7336
rect 14424 7324 14430 7336
rect 14424 7296 14469 7324
rect 14424 7284 14430 7296
rect 8113 7259 8171 7265
rect 8113 7256 8125 7259
rect 7392 7228 8125 7256
rect 7193 7219 7251 7225
rect 8113 7225 8125 7228
rect 8159 7225 8171 7259
rect 8113 7219 8171 7225
rect 9033 7259 9091 7265
rect 9033 7225 9045 7259
rect 9079 7256 9091 7259
rect 12526 7256 12532 7268
rect 9079 7228 12532 7256
rect 9079 7225 9091 7228
rect 9033 7219 9091 7225
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 3513 7191 3571 7197
rect 3513 7188 3525 7191
rect 3292 7160 3525 7188
rect 3292 7148 3298 7160
rect 3513 7157 3525 7160
rect 3559 7157 3571 7191
rect 3513 7151 3571 7157
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7188 5135 7191
rect 5258 7188 5264 7200
rect 5123 7160 5264 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 5537 7191 5595 7197
rect 5537 7157 5549 7191
rect 5583 7188 5595 7191
rect 5718 7188 5724 7200
rect 5583 7160 5724 7188
rect 5583 7157 5595 7160
rect 5537 7151 5595 7157
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 7208 7188 7236 7219
rect 12526 7216 12532 7228
rect 12584 7216 12590 7268
rect 7466 7188 7472 7200
rect 7208 7160 7472 7188
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 8938 7148 8944 7200
rect 8996 7188 9002 7200
rect 9585 7191 9643 7197
rect 9585 7188 9597 7191
rect 8996 7160 9597 7188
rect 8996 7148 9002 7160
rect 9585 7157 9597 7160
rect 9631 7157 9643 7191
rect 9585 7151 9643 7157
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 10192 7160 10425 7188
rect 10192 7148 10198 7160
rect 10413 7157 10425 7160
rect 10459 7188 10471 7191
rect 11054 7188 11060 7200
rect 10459 7160 11060 7188
rect 10459 7157 10471 7160
rect 10413 7151 10471 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 11793 7191 11851 7197
rect 11793 7188 11805 7191
rect 11204 7160 11805 7188
rect 11204 7148 11210 7160
rect 11793 7157 11805 7160
rect 11839 7188 11851 7191
rect 12066 7188 12072 7200
rect 11839 7160 12072 7188
rect 11839 7157 11851 7160
rect 11793 7151 11851 7157
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 12250 7188 12256 7200
rect 12211 7160 12256 7188
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12802 7188 12808 7200
rect 12492 7160 12808 7188
rect 12492 7148 12498 7160
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 13814 7148 13820 7200
rect 13872 7188 13878 7200
rect 14001 7191 14059 7197
rect 14001 7188 14013 7191
rect 13872 7160 14013 7188
rect 13872 7148 13878 7160
rect 14001 7157 14013 7160
rect 14047 7157 14059 7191
rect 14001 7151 14059 7157
rect 1104 7098 15732 7120
rect 1104 7046 3420 7098
rect 3472 7046 3484 7098
rect 3536 7046 3548 7098
rect 3600 7046 3612 7098
rect 3664 7046 8296 7098
rect 8348 7046 8360 7098
rect 8412 7046 8424 7098
rect 8476 7046 8488 7098
rect 8540 7046 13172 7098
rect 13224 7046 13236 7098
rect 13288 7046 13300 7098
rect 13352 7046 13364 7098
rect 13416 7046 15732 7098
rect 1104 7024 15732 7046
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 2924 6956 7880 6984
rect 2924 6944 2930 6956
rect 7852 6916 7880 6956
rect 8846 6944 8852 6996
rect 8904 6984 8910 6996
rect 10594 6984 10600 6996
rect 8904 6956 10600 6984
rect 8904 6944 8910 6956
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 10962 6984 10968 6996
rect 10923 6956 10968 6984
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 11606 6984 11612 6996
rect 11112 6956 11612 6984
rect 11112 6944 11118 6956
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 11974 6944 11980 6996
rect 12032 6984 12038 6996
rect 12342 6984 12348 6996
rect 12032 6956 12348 6984
rect 12032 6944 12038 6956
rect 12342 6944 12348 6956
rect 12400 6984 12406 6996
rect 12400 6956 12572 6984
rect 12400 6944 12406 6956
rect 12544 6925 12572 6956
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 13173 6987 13231 6993
rect 13173 6984 13185 6987
rect 12860 6956 13185 6984
rect 12860 6944 12866 6956
rect 13173 6953 13185 6956
rect 13219 6953 13231 6987
rect 13173 6947 13231 6953
rect 12529 6919 12587 6925
rect 6472 6888 7788 6916
rect 7852 6888 12480 6916
rect 2130 6848 2136 6860
rect 1872 6820 2136 6848
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 1872 6789 1900 6820
rect 2130 6808 2136 6820
rect 2188 6848 2194 6860
rect 4249 6851 4307 6857
rect 2188 6820 2452 6848
rect 2188 6808 2194 6820
rect 2424 6789 2452 6820
rect 4249 6817 4261 6851
rect 4295 6848 4307 6851
rect 4430 6848 4436 6860
rect 4295 6820 4436 6848
rect 4295 6817 4307 6820
rect 4249 6811 4307 6817
rect 4430 6808 4436 6820
rect 4488 6808 4494 6860
rect 5077 6851 5135 6857
rect 5077 6817 5089 6851
rect 5123 6848 5135 6851
rect 5258 6848 5264 6860
rect 5123 6820 5264 6848
rect 5123 6817 5135 6820
rect 5077 6811 5135 6817
rect 5258 6808 5264 6820
rect 5316 6848 5322 6860
rect 5537 6851 5595 6857
rect 5537 6848 5549 6851
rect 5316 6820 5549 6848
rect 5316 6808 5322 6820
rect 5537 6817 5549 6820
rect 5583 6817 5595 6851
rect 5537 6811 5595 6817
rect 6181 6851 6239 6857
rect 6181 6817 6193 6851
rect 6227 6817 6239 6851
rect 6472 6848 6500 6888
rect 6181 6811 6239 6817
rect 6380 6820 6500 6848
rect 6549 6851 6607 6857
rect 1857 6783 1915 6789
rect 1857 6780 1869 6783
rect 1636 6752 1869 6780
rect 1636 6740 1642 6752
rect 1857 6749 1869 6752
rect 1903 6749 1915 6783
rect 1857 6743 1915 6749
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 2409 6783 2467 6789
rect 2087 6752 2360 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 2332 6656 2360 6752
rect 2409 6749 2421 6783
rect 2455 6749 2467 6783
rect 3970 6780 3976 6792
rect 3931 6752 3976 6780
rect 2409 6743 2467 6749
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 4341 6783 4399 6789
rect 4120 6752 4165 6780
rect 4120 6740 4126 6752
rect 4341 6749 4353 6783
rect 4387 6749 4399 6783
rect 5166 6780 5172 6792
rect 5127 6752 5172 6780
rect 4341 6743 4399 6749
rect 3234 6672 3240 6724
rect 3292 6712 3298 6724
rect 4356 6712 4384 6743
rect 5166 6740 5172 6752
rect 5224 6780 5230 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 5224 6752 5457 6780
rect 5224 6740 5230 6752
rect 5445 6749 5457 6752
rect 5491 6780 5503 6783
rect 6196 6780 6224 6811
rect 5491 6752 6224 6780
rect 5491 6749 5503 6752
rect 5445 6743 5503 6749
rect 6270 6740 6276 6792
rect 6328 6780 6334 6792
rect 6380 6789 6408 6820
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 7282 6848 7288 6860
rect 6595 6820 7288 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 7282 6808 7288 6820
rect 7340 6808 7346 6860
rect 7650 6848 7656 6860
rect 7611 6820 7656 6848
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 6328 6752 6377 6780
rect 6328 6740 6334 6752
rect 6365 6749 6377 6752
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6749 6699 6783
rect 6822 6780 6828 6792
rect 6783 6752 6828 6780
rect 6641 6743 6699 6749
rect 3292 6684 4384 6712
rect 3292 6672 3298 6684
rect 1578 6604 1584 6656
rect 1636 6644 1642 6656
rect 2133 6647 2191 6653
rect 2133 6644 2145 6647
rect 1636 6616 2145 6644
rect 1636 6604 1642 6616
rect 2133 6613 2145 6616
rect 2179 6613 2191 6647
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2133 6607 2191 6613
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 3050 6604 3056 6656
rect 3108 6644 3114 6656
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 3108 6616 3801 6644
rect 3108 6604 3114 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 3789 6607 3847 6613
rect 4893 6647 4951 6653
rect 4893 6613 4905 6647
rect 4939 6644 4951 6647
rect 4982 6644 4988 6656
rect 4939 6616 4988 6644
rect 4939 6613 4951 6616
rect 4893 6607 4951 6613
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 6472 6644 6500 6743
rect 6656 6712 6684 6743
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 7558 6780 7564 6792
rect 7519 6752 7564 6780
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 7760 6789 7788 6888
rect 8297 6851 8355 6857
rect 8297 6817 8309 6851
rect 8343 6848 8355 6851
rect 10410 6848 10416 6860
rect 8343 6820 10416 6848
rect 8343 6817 8355 6820
rect 8297 6811 8355 6817
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 10980 6820 11529 6848
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 7834 6780 7840 6792
rect 7791 6752 7840 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 7984 6752 8217 6780
rect 7984 6740 7990 6752
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 8386 6780 8392 6792
rect 8347 6752 8392 6780
rect 8205 6743 8263 6749
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 8662 6740 8668 6792
rect 8720 6780 8726 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8720 6752 9137 6780
rect 8720 6740 8726 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 6730 6712 6736 6724
rect 6656 6684 6736 6712
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 9140 6712 9168 6743
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 9272 6752 9505 6780
rect 9272 6740 9278 6752
rect 9493 6749 9505 6752
rect 9539 6780 9551 6783
rect 9539 6752 9812 6780
rect 9539 6749 9551 6752
rect 9493 6743 9551 6749
rect 9585 6715 9643 6721
rect 9585 6712 9597 6715
rect 9140 6684 9597 6712
rect 9585 6681 9597 6684
rect 9631 6681 9643 6715
rect 9585 6675 9643 6681
rect 7558 6644 7564 6656
rect 6472 6616 7564 6644
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 8536 6616 8953 6644
rect 8536 6604 8542 6616
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 9784 6644 9812 6752
rect 9858 6740 9864 6792
rect 9916 6780 9922 6792
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 9916 6752 10149 6780
rect 9916 6740 9922 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10226 6672 10232 6724
rect 10284 6712 10290 6724
rect 10321 6715 10379 6721
rect 10321 6712 10333 6715
rect 10284 6684 10333 6712
rect 10284 6672 10290 6684
rect 10321 6681 10333 6684
rect 10367 6681 10379 6715
rect 10321 6675 10379 6681
rect 10505 6715 10563 6721
rect 10505 6681 10517 6715
rect 10551 6712 10563 6715
rect 10980 6712 11008 6820
rect 11517 6817 11529 6820
rect 11563 6848 11575 6851
rect 11563 6820 12388 6848
rect 11563 6817 11575 6820
rect 11517 6811 11575 6817
rect 11118 6783 11176 6789
rect 11118 6749 11130 6783
rect 11164 6780 11176 6783
rect 11609 6783 11667 6789
rect 11609 6780 11621 6783
rect 11164 6752 11621 6780
rect 11164 6749 11176 6752
rect 11118 6743 11176 6749
rect 11609 6749 11621 6752
rect 11655 6780 11667 6783
rect 12250 6780 12256 6792
rect 11655 6752 12256 6780
rect 11655 6749 11667 6752
rect 11609 6743 11667 6749
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 12360 6789 12388 6820
rect 12345 6783 12403 6789
rect 12345 6749 12357 6783
rect 12391 6749 12403 6783
rect 12345 6743 12403 6749
rect 11214 6715 11272 6721
rect 11214 6712 11226 6715
rect 10551 6684 11226 6712
rect 10551 6681 10563 6684
rect 10505 6675 10563 6681
rect 11214 6681 11226 6684
rect 11260 6681 11272 6715
rect 12452 6712 12480 6888
rect 12529 6885 12541 6919
rect 12575 6916 12587 6919
rect 12575 6888 12756 6916
rect 12575 6885 12587 6888
rect 12529 6879 12587 6885
rect 12728 6848 12756 6888
rect 12728 6820 13124 6848
rect 12621 6783 12679 6789
rect 12621 6749 12633 6783
rect 12667 6780 12679 6783
rect 12894 6780 12900 6792
rect 12667 6752 12900 6780
rect 12667 6749 12679 6752
rect 12621 6743 12679 6749
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 13096 6789 13124 6820
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 14093 6851 14151 6857
rect 14093 6848 14105 6851
rect 13780 6820 14105 6848
rect 13780 6808 13786 6820
rect 14093 6817 14105 6820
rect 14139 6817 14151 6851
rect 14366 6848 14372 6860
rect 14327 6820 14372 6848
rect 14093 6811 14151 6817
rect 14366 6808 14372 6820
rect 14424 6808 14430 6860
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 13630 6740 13636 6792
rect 13688 6780 13694 6792
rect 14384 6780 14412 6808
rect 13688 6752 14412 6780
rect 13688 6740 13694 6752
rect 12986 6712 12992 6724
rect 12452 6684 12992 6712
rect 11214 6675 11272 6681
rect 12986 6672 12992 6684
rect 13044 6672 13050 6724
rect 12069 6647 12127 6653
rect 12069 6644 12081 6647
rect 9784 6616 12081 6644
rect 8941 6607 8999 6613
rect 12069 6613 12081 6616
rect 12115 6613 12127 6647
rect 12069 6607 12127 6613
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 14642 6644 14648 6656
rect 12216 6616 14648 6644
rect 12216 6604 12222 6616
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 1104 6554 15732 6576
rect 1104 6502 5858 6554
rect 5910 6502 5922 6554
rect 5974 6502 5986 6554
rect 6038 6502 6050 6554
rect 6102 6502 10734 6554
rect 10786 6502 10798 6554
rect 10850 6502 10862 6554
rect 10914 6502 10926 6554
rect 10978 6502 15732 6554
rect 1104 6480 15732 6502
rect 1670 6400 1676 6452
rect 1728 6440 1734 6452
rect 1857 6443 1915 6449
rect 1857 6440 1869 6443
rect 1728 6412 1869 6440
rect 1728 6400 1734 6412
rect 1857 6409 1869 6412
rect 1903 6409 1915 6443
rect 1857 6403 1915 6409
rect 3973 6443 4031 6449
rect 3973 6409 3985 6443
rect 4019 6440 4031 6443
rect 4062 6440 4068 6452
rect 4019 6412 4068 6440
rect 4019 6409 4031 6412
rect 3973 6403 4031 6409
rect 1872 6304 1900 6403
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4430 6440 4436 6452
rect 4391 6412 4436 6440
rect 4430 6400 4436 6412
rect 4488 6400 4494 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 5092 6412 7941 6440
rect 3234 6332 3240 6384
rect 3292 6372 3298 6384
rect 3329 6375 3387 6381
rect 3329 6372 3341 6375
rect 3292 6344 3341 6372
rect 3292 6332 3298 6344
rect 3329 6341 3341 6344
rect 3375 6341 3387 6375
rect 3329 6335 3387 6341
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 1872 6276 2145 6304
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 1578 6196 1584 6248
rect 1636 6236 1642 6248
rect 1765 6239 1823 6245
rect 1765 6236 1777 6239
rect 1636 6208 1777 6236
rect 1636 6196 1642 6208
rect 1765 6205 1777 6208
rect 1811 6236 1823 6239
rect 2317 6239 2375 6245
rect 2317 6236 2329 6239
rect 1811 6208 2329 6236
rect 1811 6205 1823 6208
rect 1765 6199 1823 6205
rect 2317 6205 2329 6208
rect 2363 6205 2375 6239
rect 3344 6236 3372 6335
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3697 6307 3755 6313
rect 3697 6304 3709 6307
rect 3467 6276 3709 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 3697 6273 3709 6276
rect 3743 6304 3755 6307
rect 4448 6304 4476 6400
rect 4890 6372 4896 6384
rect 4632 6344 4896 6372
rect 4632 6313 4660 6344
rect 4890 6332 4896 6344
rect 4948 6372 4954 6384
rect 5092 6381 5120 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 8846 6440 8852 6452
rect 7929 6403 7987 6409
rect 8036 6412 8852 6440
rect 5077 6375 5135 6381
rect 5077 6372 5089 6375
rect 4948 6344 5089 6372
rect 4948 6332 4954 6344
rect 5077 6341 5089 6344
rect 5123 6341 5135 6375
rect 5077 6335 5135 6341
rect 6362 6332 6368 6384
rect 6420 6372 6426 6384
rect 6822 6372 6828 6384
rect 6420 6344 6828 6372
rect 6420 6332 6426 6344
rect 6822 6332 6828 6344
rect 6880 6372 6886 6384
rect 7009 6375 7067 6381
rect 7009 6372 7021 6375
rect 6880 6344 7021 6372
rect 6880 6332 6886 6344
rect 7009 6341 7021 6344
rect 7055 6341 7067 6375
rect 7009 6335 7067 6341
rect 7098 6332 7104 6384
rect 7156 6372 7162 6384
rect 8036 6372 8064 6412
rect 8846 6400 8852 6412
rect 8904 6400 8910 6452
rect 9582 6440 9588 6452
rect 9543 6412 9588 6440
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 11698 6440 11704 6452
rect 11072 6412 11704 6440
rect 11072 6384 11100 6412
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 11790 6400 11796 6452
rect 11848 6440 11854 6452
rect 14274 6440 14280 6452
rect 11848 6412 14280 6440
rect 11848 6400 11854 6412
rect 14274 6400 14280 6412
rect 14332 6400 14338 6452
rect 7156 6344 7201 6372
rect 7944 6344 8064 6372
rect 7156 6332 7162 6344
rect 3743 6276 4476 6304
rect 4617 6307 4675 6313
rect 3743 6273 3755 6276
rect 3697 6267 3755 6273
rect 4617 6273 4629 6307
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 5626 6304 5632 6316
rect 5587 6276 5632 6304
rect 4709 6267 4767 6273
rect 3789 6239 3847 6245
rect 3789 6236 3801 6239
rect 3344 6208 3801 6236
rect 2317 6199 2375 6205
rect 3789 6205 3801 6208
rect 3835 6205 3847 6239
rect 4724 6236 4752 6267
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 6270 6304 6276 6316
rect 5859 6276 6276 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6304 6975 6307
rect 7190 6304 7196 6316
rect 6963 6276 7196 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 4982 6236 4988 6248
rect 4724 6208 4988 6236
rect 3789 6199 3847 6205
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 5537 6239 5595 6245
rect 5537 6205 5549 6239
rect 5583 6236 5595 6239
rect 7944 6236 7972 6344
rect 8110 6332 8116 6384
rect 8168 6372 8174 6384
rect 8478 6372 8484 6384
rect 8168 6344 8484 6372
rect 8168 6332 8174 6344
rect 8220 6313 8248 6344
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 8570 6332 8576 6384
rect 8628 6372 8634 6384
rect 8628 6344 8892 6372
rect 8628 6332 8634 6344
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6273 8263 6307
rect 8864 6304 8892 6344
rect 9306 6332 9312 6384
rect 9364 6372 9370 6384
rect 9677 6375 9735 6381
rect 9677 6372 9689 6375
rect 9364 6344 9689 6372
rect 9364 6332 9370 6344
rect 9677 6341 9689 6344
rect 9723 6372 9735 6375
rect 10505 6375 10563 6381
rect 10505 6372 10517 6375
rect 9723 6344 10517 6372
rect 9723 6341 9735 6344
rect 9677 6335 9735 6341
rect 10505 6341 10517 6344
rect 10551 6341 10563 6375
rect 10505 6335 10563 6341
rect 10597 6375 10655 6381
rect 10597 6341 10609 6375
rect 10643 6372 10655 6375
rect 11054 6372 11060 6384
rect 10643 6344 11060 6372
rect 10643 6341 10655 6344
rect 10597 6335 10655 6341
rect 11054 6332 11060 6344
rect 11112 6332 11118 6384
rect 11330 6332 11336 6384
rect 11388 6372 11394 6384
rect 11388 6344 14136 6372
rect 11388 6332 11394 6344
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 8864 6276 9505 6304
rect 8205 6267 8263 6273
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 9950 6264 9956 6316
rect 10008 6304 10014 6316
rect 10778 6304 10784 6316
rect 10008 6276 10784 6304
rect 10008 6264 10014 6276
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 11790 6304 11796 6316
rect 11751 6276 11796 6304
rect 11790 6264 11796 6276
rect 11848 6264 11854 6316
rect 11974 6304 11980 6316
rect 11935 6276 11980 6304
rect 11974 6264 11980 6276
rect 12032 6264 12038 6316
rect 12802 6304 12808 6316
rect 12763 6276 12808 6304
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 12897 6307 12955 6313
rect 12897 6273 12909 6307
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 5583 6208 7972 6236
rect 5583 6205 5595 6208
rect 5537 6199 5595 6205
rect 8018 6196 8024 6248
rect 8076 6236 8082 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 8076 6208 8125 6236
rect 8076 6196 8082 6208
rect 8113 6205 8125 6208
rect 8159 6236 8171 6239
rect 8573 6239 8631 6245
rect 8573 6236 8585 6239
rect 8159 6208 8585 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 8573 6205 8585 6208
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 9582 6196 9588 6248
rect 9640 6236 9646 6248
rect 11146 6236 11152 6248
rect 9640 6208 11152 6236
rect 9640 6196 9646 6208
rect 11146 6196 11152 6208
rect 11204 6196 11210 6248
rect 11606 6196 11612 6248
rect 11664 6236 11670 6248
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 11664 6208 11713 6236
rect 11664 6196 11670 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 2590 6128 2596 6180
rect 2648 6168 2654 6180
rect 2648 6140 2774 6168
rect 2648 6128 2654 6140
rect 2038 6100 2044 6112
rect 1999 6072 2044 6100
rect 2038 6060 2044 6072
rect 2096 6060 2102 6112
rect 2746 6100 2774 6140
rect 3234 6128 3240 6180
rect 3292 6168 3298 6180
rect 6362 6168 6368 6180
rect 3292 6140 6368 6168
rect 3292 6128 3298 6140
rect 6362 6128 6368 6140
rect 6420 6128 6426 6180
rect 7285 6171 7343 6177
rect 7285 6137 7297 6171
rect 7331 6168 7343 6171
rect 9122 6168 9128 6180
rect 7331 6140 9128 6168
rect 7331 6137 7343 6140
rect 7285 6131 7343 6137
rect 9122 6128 9128 6140
rect 9180 6128 9186 6180
rect 9306 6168 9312 6180
rect 9267 6140 9312 6168
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 9490 6128 9496 6180
rect 9548 6168 9554 6180
rect 9861 6171 9919 6177
rect 9861 6168 9873 6171
rect 9548 6140 9873 6168
rect 9548 6128 9554 6140
rect 9861 6137 9873 6140
rect 9907 6137 9919 6171
rect 9861 6131 9919 6137
rect 10134 6128 10140 6180
rect 10192 6168 10198 6180
rect 10318 6168 10324 6180
rect 10192 6140 10324 6168
rect 10192 6128 10198 6140
rect 10318 6128 10324 6140
rect 10376 6128 10382 6180
rect 10505 6171 10563 6177
rect 10505 6137 10517 6171
rect 10551 6168 10563 6171
rect 12912 6168 12940 6267
rect 12986 6264 12992 6316
rect 13044 6304 13050 6316
rect 13127 6307 13185 6313
rect 13044 6276 13089 6304
rect 13044 6264 13050 6276
rect 13127 6273 13139 6307
rect 13173 6304 13185 6307
rect 13814 6304 13820 6316
rect 13173 6276 13820 6304
rect 13173 6273 13185 6276
rect 13127 6267 13185 6273
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 14108 6313 14136 6344
rect 14292 6313 14320 6400
rect 14093 6307 14151 6313
rect 14093 6273 14105 6307
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 13265 6239 13323 6245
rect 13265 6236 13277 6239
rect 13004 6208 13277 6236
rect 13004 6180 13032 6208
rect 13265 6205 13277 6208
rect 13311 6236 13323 6239
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13311 6208 14013 6236
rect 13311 6205 13323 6208
rect 13265 6199 13323 6205
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 14185 6239 14243 6245
rect 14185 6205 14197 6239
rect 14231 6236 14243 6239
rect 14550 6236 14556 6248
rect 14231 6208 14556 6236
rect 14231 6205 14243 6208
rect 14185 6199 14243 6205
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 10551 6140 11161 6168
rect 10551 6137 10563 6140
rect 10505 6131 10563 6137
rect 5537 6103 5595 6109
rect 5537 6100 5549 6103
rect 2746 6072 5549 6100
rect 5537 6069 5549 6072
rect 5583 6069 5595 6103
rect 5537 6063 5595 6069
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6100 5687 6103
rect 5994 6100 6000 6112
rect 5675 6072 6000 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 6733 6103 6791 6109
rect 6733 6069 6745 6103
rect 6779 6100 6791 6103
rect 7098 6100 7104 6112
rect 6779 6072 7104 6100
rect 6779 6069 6791 6072
rect 6733 6063 6791 6069
rect 7098 6060 7104 6072
rect 7156 6060 7162 6112
rect 8938 6060 8944 6112
rect 8996 6100 9002 6112
rect 10870 6100 10876 6112
rect 8996 6072 10876 6100
rect 8996 6060 9002 6072
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11133 6100 11161 6140
rect 11900 6140 12940 6168
rect 11900 6100 11928 6140
rect 12986 6128 12992 6180
rect 13044 6128 13050 6180
rect 12158 6100 12164 6112
rect 11020 6072 11065 6100
rect 11133 6072 11928 6100
rect 12119 6072 12164 6100
rect 11020 6060 11026 6072
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12250 6060 12256 6112
rect 12308 6100 12314 6112
rect 12621 6103 12679 6109
rect 12621 6100 12633 6103
rect 12308 6072 12633 6100
rect 12308 6060 12314 6072
rect 12621 6069 12633 6072
rect 12667 6069 12679 6103
rect 12621 6063 12679 6069
rect 14461 6103 14519 6109
rect 14461 6069 14473 6103
rect 14507 6100 14519 6103
rect 14826 6100 14832 6112
rect 14507 6072 14832 6100
rect 14507 6069 14519 6072
rect 14461 6063 14519 6069
rect 14826 6060 14832 6072
rect 14884 6060 14890 6112
rect 1104 6010 15732 6032
rect 1104 5958 3420 6010
rect 3472 5958 3484 6010
rect 3536 5958 3548 6010
rect 3600 5958 3612 6010
rect 3664 5958 8296 6010
rect 8348 5958 8360 6010
rect 8412 5958 8424 6010
rect 8476 5958 8488 6010
rect 8540 5958 13172 6010
rect 13224 5958 13236 6010
rect 13288 5958 13300 6010
rect 13352 5958 13364 6010
rect 13416 5958 15732 6010
rect 1104 5936 15732 5958
rect 2038 5856 2044 5908
rect 2096 5896 2102 5908
rect 8297 5899 8355 5905
rect 2096 5868 7604 5896
rect 2096 5856 2102 5868
rect 3234 5828 3240 5840
rect 3195 5800 3240 5828
rect 3234 5788 3240 5800
rect 3292 5788 3298 5840
rect 5721 5831 5779 5837
rect 5721 5828 5733 5831
rect 4448 5800 5733 5828
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5729 1915 5763
rect 3970 5760 3976 5772
rect 3883 5732 3976 5760
rect 1857 5723 1915 5729
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 1670 5652 1676 5704
rect 1728 5692 1734 5704
rect 1728 5664 1773 5692
rect 1728 5652 1734 5664
rect 1872 5624 1900 5723
rect 3970 5720 3976 5732
rect 4028 5760 4034 5772
rect 4448 5769 4476 5800
rect 5721 5797 5733 5800
rect 5767 5797 5779 5831
rect 5721 5791 5779 5797
rect 7101 5831 7159 5837
rect 7101 5797 7113 5831
rect 7147 5828 7159 5831
rect 7374 5828 7380 5840
rect 7147 5800 7380 5828
rect 7147 5797 7159 5800
rect 7101 5791 7159 5797
rect 7374 5788 7380 5800
rect 7432 5788 7438 5840
rect 7576 5828 7604 5868
rect 8297 5865 8309 5899
rect 8343 5896 8355 5899
rect 9214 5896 9220 5908
rect 8343 5868 9220 5896
rect 8343 5865 8355 5868
rect 8297 5859 8355 5865
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 11517 5899 11575 5905
rect 11517 5896 11529 5899
rect 9324 5868 11529 5896
rect 7576 5800 8524 5828
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4028 5732 4445 5760
rect 4028 5720 4034 5732
rect 4433 5729 4445 5732
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 5905 5763 5963 5769
rect 5905 5729 5917 5763
rect 5951 5760 5963 5763
rect 6365 5763 6423 5769
rect 6365 5760 6377 5763
rect 5951 5732 6377 5760
rect 5951 5729 5963 5732
rect 5905 5723 5963 5729
rect 6365 5729 6377 5732
rect 6411 5760 6423 5763
rect 6411 5732 6960 5760
rect 6411 5729 6423 5732
rect 6365 5723 6423 5729
rect 6932 5704 6960 5732
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5692 2007 5695
rect 2130 5692 2136 5704
rect 1995 5664 2136 5692
rect 1995 5661 2007 5664
rect 1949 5655 2007 5661
rect 2130 5652 2136 5664
rect 2188 5652 2194 5704
rect 2406 5692 2412 5704
rect 2367 5664 2412 5692
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5692 3111 5695
rect 3099 5664 4016 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 2314 5624 2320 5636
rect 1872 5596 2320 5624
rect 2314 5584 2320 5596
rect 2372 5624 2378 5636
rect 3988 5624 4016 5664
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4341 5695 4399 5701
rect 4341 5692 4353 5695
rect 4120 5664 4353 5692
rect 4120 5652 4126 5664
rect 4341 5661 4353 5664
rect 4387 5661 4399 5695
rect 4341 5655 4399 5661
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5692 5319 5695
rect 5350 5692 5356 5704
rect 5307 5664 5356 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 5994 5652 6000 5704
rect 6052 5692 6058 5704
rect 6273 5695 6331 5701
rect 6273 5692 6285 5695
rect 6052 5664 6285 5692
rect 6052 5652 6058 5664
rect 6273 5661 6285 5664
rect 6319 5692 6331 5695
rect 6825 5695 6883 5701
rect 6825 5692 6837 5695
rect 6319 5664 6837 5692
rect 6319 5661 6331 5664
rect 6273 5655 6331 5661
rect 6825 5661 6837 5664
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 8018 5692 8024 5704
rect 6972 5664 7065 5692
rect 7931 5664 8024 5692
rect 6972 5652 6978 5664
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 8110 5652 8116 5704
rect 8168 5692 8174 5704
rect 8386 5692 8392 5704
rect 8168 5664 8213 5692
rect 8347 5664 8392 5692
rect 8168 5652 8174 5664
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 8496 5692 8524 5800
rect 9324 5769 9352 5868
rect 11517 5865 11529 5868
rect 11563 5865 11575 5899
rect 11517 5859 11575 5865
rect 9493 5831 9551 5837
rect 9493 5797 9505 5831
rect 9539 5828 9551 5831
rect 9858 5828 9864 5840
rect 9539 5800 9864 5828
rect 9539 5797 9551 5800
rect 9493 5791 9551 5797
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 10042 5828 10048 5840
rect 10003 5800 10048 5828
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 10965 5831 11023 5837
rect 10965 5828 10977 5831
rect 10152 5800 10977 5828
rect 9309 5763 9367 5769
rect 9309 5729 9321 5763
rect 9355 5729 9367 5763
rect 10152 5760 10180 5800
rect 10965 5797 10977 5800
rect 11011 5797 11023 5831
rect 11532 5828 11560 5859
rect 12802 5856 12808 5908
rect 12860 5896 12866 5908
rect 13449 5899 13507 5905
rect 13449 5896 13461 5899
rect 12860 5868 13461 5896
rect 12860 5856 12866 5868
rect 13449 5865 13461 5868
rect 13495 5865 13507 5899
rect 13449 5859 13507 5865
rect 14458 5856 14464 5908
rect 14516 5896 14522 5908
rect 14829 5899 14887 5905
rect 14829 5896 14841 5899
rect 14516 5868 14841 5896
rect 14516 5856 14522 5868
rect 14829 5865 14841 5868
rect 14875 5865 14887 5899
rect 14829 5859 14887 5865
rect 11974 5828 11980 5840
rect 11532 5800 11980 5828
rect 10965 5791 11023 5797
rect 9309 5723 9367 5729
rect 9600 5732 10180 5760
rect 10980 5760 11008 5791
rect 11974 5788 11980 5800
rect 12032 5828 12038 5840
rect 12032 5800 12112 5828
rect 12032 5788 12038 5800
rect 10980 5732 11652 5760
rect 9600 5701 9628 5732
rect 9585 5695 9643 5701
rect 8496 5664 9444 5692
rect 6730 5624 6736 5636
rect 2372 5596 3832 5624
rect 3988 5596 6736 5624
rect 2372 5584 2378 5596
rect 1397 5559 1455 5565
rect 1397 5525 1409 5559
rect 1443 5556 1455 5559
rect 1578 5556 1584 5568
rect 1443 5528 1584 5556
rect 1443 5525 1455 5528
rect 1397 5519 1455 5525
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 2590 5556 2596 5568
rect 2551 5528 2596 5556
rect 2590 5516 2596 5528
rect 2648 5516 2654 5568
rect 3804 5565 3832 5596
rect 6730 5584 6736 5596
rect 6788 5584 6794 5636
rect 7098 5624 7104 5636
rect 7059 5596 7104 5624
rect 7098 5584 7104 5596
rect 7156 5584 7162 5636
rect 8036 5624 8064 5652
rect 9309 5627 9367 5633
rect 9309 5624 9321 5627
rect 8036 5596 9321 5624
rect 9309 5593 9321 5596
rect 9355 5593 9367 5627
rect 9416 5624 9444 5664
rect 9585 5661 9597 5695
rect 9631 5661 9643 5695
rect 9585 5655 9643 5661
rect 10330 5695 10388 5701
rect 10330 5661 10342 5695
rect 10376 5691 10388 5695
rect 10594 5692 10600 5704
rect 10428 5691 10600 5692
rect 10376 5664 10600 5691
rect 10376 5663 10456 5664
rect 10376 5661 10388 5663
rect 10330 5655 10388 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 10778 5692 10784 5704
rect 10739 5664 10784 5692
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 10962 5692 10968 5704
rect 10923 5664 10968 5692
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 11624 5701 11652 5732
rect 12084 5701 12112 5800
rect 13998 5788 14004 5840
rect 14056 5828 14062 5840
rect 14274 5828 14280 5840
rect 14056 5800 14280 5828
rect 14056 5788 14062 5800
rect 14274 5788 14280 5800
rect 14332 5828 14338 5840
rect 14332 5800 14688 5828
rect 14332 5788 14338 5800
rect 14366 5760 14372 5772
rect 14327 5732 14372 5760
rect 14366 5720 14372 5732
rect 14424 5720 14430 5772
rect 14461 5763 14519 5769
rect 14461 5729 14473 5763
rect 14507 5760 14519 5763
rect 14550 5760 14556 5772
rect 14507 5732 14556 5760
rect 14507 5729 14519 5732
rect 14461 5723 14519 5729
rect 14550 5720 14556 5732
rect 14608 5720 14614 5772
rect 11425 5695 11483 5701
rect 11425 5661 11437 5695
rect 11471 5661 11483 5695
rect 11425 5655 11483 5661
rect 11609 5695 11667 5701
rect 11609 5661 11621 5695
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5692 12311 5695
rect 12342 5692 12348 5704
rect 12299 5664 12348 5692
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 9766 5624 9772 5636
rect 9416 5596 9772 5624
rect 9309 5587 9367 5593
rect 9766 5584 9772 5596
rect 9824 5584 9830 5636
rect 10045 5627 10103 5633
rect 10045 5593 10057 5627
rect 10091 5624 10103 5627
rect 10091 5596 10364 5624
rect 10091 5593 10103 5596
rect 10045 5587 10103 5593
rect 10336 5568 10364 5596
rect 10502 5584 10508 5636
rect 10560 5624 10566 5636
rect 11440 5624 11468 5655
rect 12342 5652 12348 5664
rect 12400 5652 12406 5704
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 12897 5695 12955 5701
rect 12897 5692 12909 5695
rect 12860 5664 12909 5692
rect 12860 5652 12866 5664
rect 12897 5661 12909 5664
rect 12943 5692 12955 5695
rect 13446 5692 13452 5704
rect 12943 5664 13452 5692
rect 12943 5661 12955 5664
rect 12897 5655 12955 5661
rect 13446 5652 13452 5664
rect 13504 5652 13510 5704
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 13814 5692 13820 5704
rect 13587 5664 13820 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 13814 5652 13820 5664
rect 13872 5652 13878 5704
rect 14660 5701 14688 5800
rect 14645 5695 14703 5701
rect 14645 5661 14657 5695
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 10560 5596 11468 5624
rect 10560 5584 10566 5596
rect 14550 5584 14556 5636
rect 14608 5624 14614 5636
rect 14826 5624 14832 5636
rect 14608 5596 14832 5624
rect 14608 5584 14614 5596
rect 14826 5584 14832 5596
rect 14884 5584 14890 5636
rect 14918 5584 14924 5636
rect 14976 5584 14982 5636
rect 3789 5559 3847 5565
rect 3789 5525 3801 5559
rect 3835 5525 3847 5559
rect 3789 5519 3847 5525
rect 5169 5559 5227 5565
rect 5169 5525 5181 5559
rect 5215 5556 5227 5559
rect 5626 5556 5632 5568
rect 5215 5528 5632 5556
rect 5215 5525 5227 5528
rect 5169 5519 5227 5525
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 7834 5556 7840 5568
rect 7795 5528 7840 5556
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 9674 5556 9680 5568
rect 8260 5528 9680 5556
rect 8260 5516 8266 5528
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 10134 5516 10140 5568
rect 10192 5556 10198 5568
rect 10229 5559 10287 5565
rect 10229 5556 10241 5559
rect 10192 5528 10241 5556
rect 10192 5516 10198 5528
rect 10229 5525 10241 5528
rect 10275 5525 10287 5559
rect 10229 5519 10287 5525
rect 10318 5516 10324 5568
rect 10376 5516 10382 5568
rect 11790 5516 11796 5568
rect 11848 5556 11854 5568
rect 12161 5559 12219 5565
rect 12161 5556 12173 5559
rect 11848 5528 12173 5556
rect 11848 5516 11854 5528
rect 12161 5525 12173 5528
rect 12207 5525 12219 5559
rect 12802 5556 12808 5568
rect 12763 5528 12808 5556
rect 12161 5519 12219 5525
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 13998 5516 14004 5568
rect 14056 5556 14062 5568
rect 14936 5556 14964 5584
rect 14056 5528 14964 5556
rect 14056 5516 14062 5528
rect 1104 5466 15732 5488
rect 1104 5414 5858 5466
rect 5910 5414 5922 5466
rect 5974 5414 5986 5466
rect 6038 5414 6050 5466
rect 6102 5414 10734 5466
rect 10786 5414 10798 5466
rect 10850 5414 10862 5466
rect 10914 5414 10926 5466
rect 10978 5414 15732 5466
rect 1104 5392 15732 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5321 1639 5355
rect 1581 5315 1639 5321
rect 2593 5355 2651 5361
rect 2593 5321 2605 5355
rect 2639 5352 2651 5355
rect 2866 5352 2872 5364
rect 2639 5324 2872 5352
rect 2639 5321 2651 5324
rect 2593 5315 2651 5321
rect 1596 5284 1624 5315
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 3142 5312 3148 5364
rect 3200 5352 3206 5364
rect 3200 5324 6868 5352
rect 3200 5312 3206 5324
rect 4614 5284 4620 5296
rect 1596 5256 4620 5284
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 6840 5284 6868 5324
rect 6914 5312 6920 5364
rect 6972 5352 6978 5364
rect 7009 5355 7067 5361
rect 7009 5352 7021 5355
rect 6972 5324 7021 5352
rect 6972 5312 6978 5324
rect 7009 5321 7021 5324
rect 7055 5321 7067 5355
rect 9766 5352 9772 5364
rect 7009 5315 7067 5321
rect 8956 5324 9772 5352
rect 8956 5284 8984 5324
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 10502 5352 10508 5364
rect 9916 5324 10508 5352
rect 9916 5312 9922 5324
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 11606 5352 11612 5364
rect 11567 5324 11612 5352
rect 11606 5312 11612 5324
rect 11664 5312 11670 5364
rect 12986 5312 12992 5364
rect 13044 5352 13050 5364
rect 13173 5355 13231 5361
rect 13173 5352 13185 5355
rect 13044 5324 13185 5352
rect 13044 5312 13050 5324
rect 13173 5321 13185 5324
rect 13219 5321 13231 5355
rect 14182 5352 14188 5364
rect 14143 5324 14188 5352
rect 13173 5315 13231 5321
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 11514 5284 11520 5296
rect 6840 5256 8984 5284
rect 9692 5256 11520 5284
rect 1394 5216 1400 5228
rect 1355 5188 1400 5216
rect 1394 5176 1400 5188
rect 1452 5176 1458 5228
rect 2406 5216 2412 5228
rect 2367 5188 2412 5216
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5216 3111 5219
rect 3142 5216 3148 5228
rect 3099 5188 3148 5216
rect 3099 5185 3111 5188
rect 3053 5179 3111 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5185 3939 5219
rect 3881 5179 3939 5185
rect 3896 5148 3924 5179
rect 3970 5176 3976 5228
rect 4028 5216 4034 5228
rect 4249 5219 4307 5225
rect 4028 5188 4073 5216
rect 4028 5176 4034 5188
rect 4249 5185 4261 5219
rect 4295 5216 4307 5219
rect 4338 5216 4344 5228
rect 4295 5188 4344 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 4338 5176 4344 5188
rect 4396 5216 4402 5228
rect 4709 5219 4767 5225
rect 4709 5216 4721 5219
rect 4396 5188 4721 5216
rect 4396 5176 4402 5188
rect 4709 5185 4721 5188
rect 4755 5185 4767 5219
rect 4890 5216 4896 5228
rect 4851 5188 4896 5216
rect 4709 5179 4767 5185
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 4982 5176 4988 5228
rect 5040 5216 5046 5228
rect 5258 5216 5264 5228
rect 5040 5188 5085 5216
rect 5219 5188 5264 5216
rect 5040 5176 5046 5188
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5216 6975 5219
rect 7006 5216 7012 5228
rect 6963 5188 7012 5216
rect 6963 5185 6975 5188
rect 6917 5179 6975 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 7101 5219 7159 5225
rect 7101 5185 7113 5219
rect 7147 5216 7159 5219
rect 7745 5219 7803 5225
rect 7745 5216 7757 5219
rect 7147 5188 7757 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7745 5185 7757 5188
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 7929 5219 7987 5225
rect 7929 5185 7941 5219
rect 7975 5185 7987 5219
rect 7929 5179 7987 5185
rect 5166 5148 5172 5160
rect 3896 5120 4292 5148
rect 5127 5120 5172 5148
rect 4264 5092 4292 5120
rect 5166 5108 5172 5120
rect 5224 5108 5230 5160
rect 6546 5108 6552 5160
rect 6604 5148 6610 5160
rect 7944 5148 7972 5179
rect 8018 5176 8024 5228
rect 8076 5216 8082 5228
rect 8297 5219 8355 5225
rect 8076 5188 8248 5216
rect 8076 5176 8082 5188
rect 6604 5120 7972 5148
rect 8220 5148 8248 5188
rect 8297 5185 8309 5219
rect 8343 5216 8355 5219
rect 8754 5216 8760 5228
rect 8343 5188 8760 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 8754 5176 8760 5188
rect 8812 5176 8818 5228
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 9033 5219 9091 5225
rect 9033 5216 9045 5219
rect 8996 5188 9045 5216
rect 8996 5176 9002 5188
rect 9033 5185 9045 5188
rect 9079 5185 9091 5219
rect 9033 5179 9091 5185
rect 9122 5176 9128 5228
rect 9180 5216 9186 5228
rect 9398 5216 9404 5228
rect 9180 5188 9404 5216
rect 9180 5176 9186 5188
rect 9398 5176 9404 5188
rect 9456 5176 9462 5228
rect 9692 5148 9720 5256
rect 11514 5244 11520 5256
rect 11572 5244 11578 5296
rect 13906 5244 13912 5296
rect 13964 5284 13970 5296
rect 14829 5287 14887 5293
rect 14829 5284 14841 5287
rect 13964 5256 14841 5284
rect 13964 5244 13970 5256
rect 14829 5253 14841 5256
rect 14875 5253 14887 5287
rect 14829 5247 14887 5253
rect 10042 5216 10048 5228
rect 10003 5188 10048 5216
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10192 5188 10237 5216
rect 10192 5176 10198 5188
rect 10318 5176 10324 5228
rect 10376 5216 10382 5228
rect 10376 5188 10421 5216
rect 10376 5176 10382 5188
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 11974 5216 11980 5228
rect 11848 5188 11893 5216
rect 11935 5188 11980 5216
rect 11848 5176 11854 5188
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5216 12127 5219
rect 12158 5216 12164 5228
rect 12115 5188 12164 5216
rect 12115 5185 12127 5188
rect 12069 5179 12127 5185
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 12805 5219 12863 5225
rect 12805 5216 12817 5219
rect 12492 5188 12817 5216
rect 12492 5176 12498 5188
rect 12805 5185 12817 5188
rect 12851 5185 12863 5219
rect 12986 5216 12992 5228
rect 12947 5188 12992 5216
rect 12805 5179 12863 5185
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 13446 5176 13452 5228
rect 13504 5216 13510 5228
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 13504 5188 14105 5216
rect 13504 5176 13510 5188
rect 14093 5185 14105 5188
rect 14139 5185 14151 5219
rect 14274 5216 14280 5228
rect 14235 5188 14280 5216
rect 14093 5179 14151 5185
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 15010 5216 15016 5228
rect 14971 5188 15016 5216
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 8220 5120 9720 5148
rect 10229 5151 10287 5157
rect 6604 5108 6610 5120
rect 10229 5117 10241 5151
rect 10275 5148 10287 5151
rect 10594 5148 10600 5160
rect 10275 5120 10600 5148
rect 10275 5117 10287 5120
rect 10229 5111 10287 5117
rect 10594 5108 10600 5120
rect 10652 5148 10658 5160
rect 11514 5148 11520 5160
rect 10652 5120 11520 5148
rect 10652 5108 10658 5120
rect 11514 5108 11520 5120
rect 11572 5148 11578 5160
rect 11885 5151 11943 5157
rect 11885 5148 11897 5151
rect 11572 5120 11897 5148
rect 11572 5108 11578 5120
rect 11885 5117 11897 5120
rect 11931 5148 11943 5151
rect 13630 5148 13636 5160
rect 11931 5120 13636 5148
rect 11931 5117 11943 5120
rect 11885 5111 11943 5117
rect 13630 5108 13636 5120
rect 13688 5108 13694 5160
rect 3145 5083 3203 5089
rect 3145 5049 3157 5083
rect 3191 5080 3203 5083
rect 4062 5080 4068 5092
rect 3191 5052 4068 5080
rect 3191 5049 3203 5052
rect 3145 5043 3203 5049
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 4246 5040 4252 5092
rect 4304 5040 4310 5092
rect 7558 5040 7564 5092
rect 7616 5080 7622 5092
rect 8110 5080 8116 5092
rect 7616 5052 8116 5080
rect 7616 5040 7622 5052
rect 8110 5040 8116 5052
rect 8168 5080 8174 5092
rect 8849 5083 8907 5089
rect 8849 5080 8861 5083
rect 8168 5052 8861 5080
rect 8168 5040 8174 5052
rect 8849 5049 8861 5052
rect 8895 5049 8907 5083
rect 8849 5043 8907 5049
rect 8938 5040 8944 5092
rect 8996 5080 9002 5092
rect 9398 5080 9404 5092
rect 8996 5052 9404 5080
rect 8996 5040 9002 5052
rect 9398 5040 9404 5052
rect 9456 5040 9462 5092
rect 10410 5040 10416 5092
rect 10468 5080 10474 5092
rect 14458 5080 14464 5092
rect 10468 5052 14464 5080
rect 10468 5040 10474 5052
rect 14458 5040 14464 5052
rect 14516 5040 14522 5092
rect 3697 5015 3755 5021
rect 3697 4981 3709 5015
rect 3743 5012 3755 5015
rect 3786 5012 3792 5024
rect 3743 4984 3792 5012
rect 3743 4981 3755 4984
rect 3697 4975 3755 4981
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 4157 5015 4215 5021
rect 4157 4981 4169 5015
rect 4203 5012 4215 5015
rect 4706 5012 4712 5024
rect 4203 4984 4712 5012
rect 4203 4981 4215 4984
rect 4157 4975 4215 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 8205 5015 8263 5021
rect 8205 4981 8217 5015
rect 8251 5012 8263 5015
rect 9122 5012 9128 5024
rect 8251 4984 9128 5012
rect 8251 4981 8263 4984
rect 8205 4975 8263 4981
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9306 5012 9312 5024
rect 9267 4984 9312 5012
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 14182 5012 14188 5024
rect 12492 4984 14188 5012
rect 12492 4972 12498 4984
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 1104 4922 15732 4944
rect 1104 4870 3420 4922
rect 3472 4870 3484 4922
rect 3536 4870 3548 4922
rect 3600 4870 3612 4922
rect 3664 4870 8296 4922
rect 8348 4870 8360 4922
rect 8412 4870 8424 4922
rect 8476 4870 8488 4922
rect 8540 4870 13172 4922
rect 13224 4870 13236 4922
rect 13288 4870 13300 4922
rect 13352 4870 13364 4922
rect 13416 4870 15732 4922
rect 1104 4848 15732 4870
rect 1673 4811 1731 4817
rect 1673 4777 1685 4811
rect 1719 4808 1731 4811
rect 1719 4780 3556 4808
rect 1719 4777 1731 4780
rect 1673 4771 1731 4777
rect 2038 4740 2044 4752
rect 1951 4712 2044 4740
rect 1964 4681 1992 4712
rect 2038 4700 2044 4712
rect 2096 4740 2102 4752
rect 2685 4743 2743 4749
rect 2685 4740 2697 4743
rect 2096 4712 2697 4740
rect 2096 4700 2102 4712
rect 2685 4709 2697 4712
rect 2731 4709 2743 4743
rect 2685 4703 2743 4709
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1949 4675 2007 4681
rect 1949 4672 1961 4675
rect 1443 4644 1961 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1949 4641 1961 4644
rect 1995 4641 2007 4675
rect 3528 4672 3556 4780
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 4028 4780 4169 4808
rect 4028 4768 4034 4780
rect 4157 4777 4169 4780
rect 4203 4777 4215 4811
rect 4157 4771 4215 4777
rect 8018 4768 8024 4820
rect 8076 4808 8082 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 8076 4780 8217 4808
rect 8076 4768 8082 4780
rect 8205 4777 8217 4780
rect 8251 4777 8263 4811
rect 8205 4771 8263 4777
rect 10229 4811 10287 4817
rect 10229 4777 10241 4811
rect 10275 4808 10287 4811
rect 10318 4808 10324 4820
rect 10275 4780 10324 4808
rect 10275 4777 10287 4780
rect 10229 4771 10287 4777
rect 10318 4768 10324 4780
rect 10376 4768 10382 4820
rect 11054 4768 11060 4820
rect 11112 4808 11118 4820
rect 12986 4808 12992 4820
rect 11112 4780 12992 4808
rect 11112 4768 11118 4780
rect 12986 4768 12992 4780
rect 13044 4768 13050 4820
rect 4062 4700 4068 4752
rect 4120 4740 4126 4752
rect 6270 4740 6276 4752
rect 4120 4712 6276 4740
rect 4120 4700 4126 4712
rect 6270 4700 6276 4712
rect 6328 4700 6334 4752
rect 8846 4700 8852 4752
rect 8904 4740 8910 4752
rect 8904 4712 11192 4740
rect 8904 4700 8910 4712
rect 4154 4672 4160 4684
rect 1949 4635 2007 4641
rect 2516 4644 3096 4672
rect 3528 4644 4160 4672
rect 1578 4604 1584 4616
rect 1539 4576 1584 4604
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 2406 4564 2412 4616
rect 2464 4604 2470 4616
rect 2516 4613 2544 4644
rect 3068 4616 3096 4644
rect 4154 4632 4160 4644
rect 4212 4632 4218 4684
rect 4338 4672 4344 4684
rect 4299 4644 4344 4672
rect 4338 4632 4344 4644
rect 4396 4672 4402 4684
rect 4801 4675 4859 4681
rect 4801 4672 4813 4675
rect 4396 4644 4813 4672
rect 4396 4632 4402 4644
rect 4801 4641 4813 4644
rect 4847 4641 4859 4675
rect 5813 4675 5871 4681
rect 5813 4672 5825 4675
rect 4801 4635 4859 4641
rect 5552 4644 5825 4672
rect 2501 4607 2559 4613
rect 2501 4604 2513 4607
rect 2464 4576 2513 4604
rect 2464 4564 2470 4576
rect 2501 4573 2513 4576
rect 2547 4573 2559 4607
rect 2501 4567 2559 4573
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4573 2651 4607
rect 3050 4604 3056 4616
rect 3011 4576 3056 4604
rect 2593 4567 2651 4573
rect 1596 4536 1624 4564
rect 1857 4539 1915 4545
rect 1857 4536 1869 4539
rect 1596 4508 1869 4536
rect 1857 4505 1869 4508
rect 1903 4536 1915 4539
rect 2130 4536 2136 4548
rect 1903 4508 2136 4536
rect 1903 4505 1915 4508
rect 1857 4499 1915 4505
rect 2130 4496 2136 4508
rect 2188 4496 2194 4548
rect 2608 4468 2636 4567
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4706 4604 4712 4616
rect 4479 4576 4712 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 5552 4613 5580 4644
rect 5813 4641 5825 4644
rect 5859 4672 5871 4675
rect 6457 4675 6515 4681
rect 6457 4672 6469 4675
rect 5859 4644 6469 4672
rect 5859 4641 5871 4644
rect 5813 4635 5871 4641
rect 6457 4641 6469 4644
rect 6503 4641 6515 4675
rect 6457 4635 6515 4641
rect 7006 4632 7012 4684
rect 7064 4672 7070 4684
rect 7285 4675 7343 4681
rect 7285 4672 7297 4675
rect 7064 4644 7297 4672
rect 7064 4632 7070 4644
rect 7285 4641 7297 4644
rect 7331 4672 7343 4675
rect 7745 4675 7803 4681
rect 7745 4672 7757 4675
rect 7331 4644 7757 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 7745 4641 7757 4644
rect 7791 4672 7803 4675
rect 7834 4672 7840 4684
rect 7791 4644 7840 4672
rect 7791 4641 7803 4644
rect 7745 4635 7803 4641
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 8662 4632 8668 4684
rect 8720 4672 8726 4684
rect 9518 4681 9546 4712
rect 9401 4675 9459 4681
rect 9401 4672 9413 4675
rect 8720 4644 9413 4672
rect 8720 4632 8726 4644
rect 9401 4641 9413 4644
rect 9447 4641 9459 4675
rect 9401 4635 9459 4641
rect 9493 4675 9551 4681
rect 9493 4641 9505 4675
rect 9539 4641 9551 4675
rect 9493 4635 9551 4641
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 10502 4672 10508 4684
rect 9732 4644 10508 4672
rect 9732 4632 9738 4644
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 5460 4536 5488 4567
rect 5718 4564 5724 4616
rect 5776 4604 5782 4616
rect 6362 4604 6368 4616
rect 5776 4576 6368 4604
rect 5776 4564 5782 4576
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 6546 4604 6552 4616
rect 6507 4576 6552 4604
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 7374 4604 7380 4616
rect 7335 4576 7380 4604
rect 7374 4564 7380 4576
rect 7432 4604 7438 4616
rect 7653 4607 7711 4613
rect 7653 4604 7665 4607
rect 7432 4576 7665 4604
rect 7432 4564 7438 4576
rect 7653 4573 7665 4576
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 8389 4607 8447 4613
rect 8389 4604 8401 4607
rect 8168 4576 8401 4604
rect 8168 4564 8174 4576
rect 8389 4573 8401 4576
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 9214 4564 9220 4616
rect 9272 4604 9278 4616
rect 9309 4607 9367 4613
rect 9309 4604 9321 4607
rect 9272 4576 9321 4604
rect 9272 4564 9278 4576
rect 9309 4573 9321 4576
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 10597 4607 10655 4613
rect 9640 4576 9685 4604
rect 9640 4564 9646 4576
rect 10597 4573 10609 4607
rect 10643 4604 10655 4607
rect 11054 4604 11060 4616
rect 10643 4576 11060 4604
rect 10643 4573 10655 4576
rect 10597 4567 10655 4573
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 5905 4539 5963 4545
rect 5905 4536 5917 4539
rect 5460 4508 5917 4536
rect 5905 4505 5917 4508
rect 5951 4536 5963 4539
rect 8938 4536 8944 4548
rect 5951 4508 8944 4536
rect 5951 4505 5963 4508
rect 5905 4499 5963 4505
rect 8938 4496 8944 4508
rect 8996 4496 9002 4548
rect 9674 4496 9680 4548
rect 9732 4536 9738 4548
rect 10226 4536 10232 4548
rect 9732 4508 10232 4536
rect 9732 4496 9738 4508
rect 10226 4496 10232 4508
rect 10284 4536 10290 4548
rect 10413 4539 10471 4545
rect 10413 4536 10425 4539
rect 10284 4508 10425 4536
rect 10284 4496 10290 4508
rect 10413 4505 10425 4508
rect 10459 4505 10471 4539
rect 11164 4536 11192 4712
rect 11882 4700 11888 4752
rect 11940 4700 11946 4752
rect 12526 4700 12532 4752
rect 12584 4740 12590 4752
rect 12584 4712 13400 4740
rect 12584 4700 12590 4712
rect 11790 4672 11796 4684
rect 11440 4644 11796 4672
rect 11440 4613 11468 4644
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 11900 4672 11928 4700
rect 11900 4644 12572 4672
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4573 11483 4607
rect 11425 4567 11483 4573
rect 11514 4564 11520 4616
rect 11572 4604 11578 4616
rect 11572 4576 11617 4604
rect 11572 4564 11578 4576
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 12544 4604 12572 4644
rect 12710 4632 12716 4684
rect 12768 4672 12774 4684
rect 12897 4675 12955 4681
rect 12897 4672 12909 4675
rect 12768 4644 12909 4672
rect 12768 4632 12774 4644
rect 12897 4641 12909 4644
rect 12943 4641 12955 4675
rect 12897 4635 12955 4641
rect 13372 4616 13400 4712
rect 14182 4700 14188 4752
rect 14240 4740 14246 4752
rect 14240 4712 14596 4740
rect 14240 4700 14246 4712
rect 14458 4672 14464 4684
rect 14419 4644 14464 4672
rect 13078 4604 13084 4616
rect 11940 4576 11985 4604
rect 12544 4576 13084 4604
rect 11940 4564 11946 4576
rect 13078 4564 13084 4576
rect 13136 4564 13142 4616
rect 13262 4604 13268 4616
rect 13223 4576 13268 4604
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 13354 4564 13360 4616
rect 13412 4613 13418 4616
rect 13412 4607 13441 4613
rect 13429 4604 13441 4607
rect 13429 4576 13505 4604
rect 13538 4584 13544 4636
rect 13596 4584 13602 4636
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 14568 4672 14596 4712
rect 14642 4700 14648 4752
rect 14700 4740 14706 4752
rect 14700 4712 14872 4740
rect 14700 4700 14706 4712
rect 14568 4644 14688 4672
rect 13429 4573 13441 4576
rect 13412 4567 13441 4573
rect 13541 4573 13553 4584
rect 13587 4573 13599 4584
rect 13541 4567 13599 4573
rect 13412 4564 13418 4567
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 13780 4576 14289 4604
rect 13780 4564 13786 4576
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14550 4604 14556 4616
rect 14463 4576 14556 4604
rect 14277 4567 14335 4573
rect 14550 4564 14556 4576
rect 14608 4564 14614 4616
rect 14660 4613 14688 4644
rect 14645 4607 14703 4613
rect 14645 4573 14657 4607
rect 14691 4573 14703 4607
rect 14645 4567 14703 4573
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4604 14795 4607
rect 14844 4604 14872 4712
rect 14783 4576 14872 4604
rect 14783 4573 14795 4576
rect 14737 4567 14795 4573
rect 11606 4536 11612 4548
rect 11164 4508 11468 4536
rect 11567 4508 11612 4536
rect 10413 4499 10471 4505
rect 2958 4468 2964 4480
rect 2608 4440 2964 4468
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 4338 4428 4344 4480
rect 4396 4468 4402 4480
rect 5261 4471 5319 4477
rect 5261 4468 5273 4471
rect 4396 4440 5273 4468
rect 4396 4428 4402 4440
rect 5261 4437 5273 4440
rect 5307 4437 5319 4471
rect 7098 4468 7104 4480
rect 7059 4440 7104 4468
rect 5261 4431 5319 4437
rect 7098 4428 7104 4440
rect 7156 4428 7162 4480
rect 8202 4428 8208 4480
rect 8260 4468 8266 4480
rect 9398 4468 9404 4480
rect 8260 4440 9404 4468
rect 8260 4428 8266 4440
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 9769 4471 9827 4477
rect 9769 4437 9781 4471
rect 9815 4468 9827 4471
rect 10134 4468 10140 4480
rect 9815 4440 10140 4468
rect 9815 4437 9827 4440
rect 9769 4431 9827 4437
rect 10134 4428 10140 4440
rect 10192 4428 10198 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11241 4471 11299 4477
rect 11241 4468 11253 4471
rect 11112 4440 11253 4468
rect 11112 4428 11118 4440
rect 11241 4437 11253 4440
rect 11287 4437 11299 4471
rect 11440 4468 11468 4508
rect 11606 4496 11612 4508
rect 11664 4496 11670 4548
rect 11747 4539 11805 4545
rect 11747 4505 11759 4539
rect 11793 4536 11805 4539
rect 12802 4536 12808 4548
rect 11793 4508 12808 4536
rect 11793 4505 11805 4508
rect 11747 4499 11805 4505
rect 12802 4496 12808 4508
rect 12860 4496 12866 4548
rect 13173 4539 13231 4545
rect 13173 4536 13185 4539
rect 12912 4508 13185 4536
rect 12526 4468 12532 4480
rect 11440 4440 12532 4468
rect 11241 4431 11299 4437
rect 12526 4428 12532 4440
rect 12584 4468 12590 4480
rect 12912 4468 12940 4508
rect 13173 4505 13185 4508
rect 13219 4505 13231 4539
rect 13173 4499 13231 4505
rect 13906 4496 13912 4548
rect 13964 4536 13970 4548
rect 14568 4536 14596 4564
rect 13964 4508 14596 4536
rect 13964 4496 13970 4508
rect 12584 4440 12940 4468
rect 12584 4428 12590 4440
rect 13078 4428 13084 4480
rect 13136 4468 13142 4480
rect 14921 4471 14979 4477
rect 14921 4468 14933 4471
rect 13136 4440 14933 4468
rect 13136 4428 13142 4440
rect 14921 4437 14933 4440
rect 14967 4437 14979 4471
rect 14921 4431 14979 4437
rect 1104 4378 15732 4400
rect 1104 4326 5858 4378
rect 5910 4326 5922 4378
rect 5974 4326 5986 4378
rect 6038 4326 6050 4378
rect 6102 4326 10734 4378
rect 10786 4326 10798 4378
rect 10850 4326 10862 4378
rect 10914 4326 10926 4378
rect 10978 4326 15732 4378
rect 1104 4304 15732 4326
rect 2958 4224 2964 4276
rect 3016 4264 3022 4276
rect 3697 4267 3755 4273
rect 3697 4264 3709 4267
rect 3016 4236 3709 4264
rect 3016 4224 3022 4236
rect 3697 4233 3709 4236
rect 3743 4233 3755 4267
rect 3697 4227 3755 4233
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 5169 4267 5227 4273
rect 5169 4264 5181 4267
rect 4764 4236 5181 4264
rect 4764 4224 4770 4236
rect 5169 4233 5181 4236
rect 5215 4233 5227 4267
rect 5169 4227 5227 4233
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 6457 4267 6515 4273
rect 6457 4264 6469 4267
rect 6420 4236 6469 4264
rect 6420 4224 6426 4236
rect 6457 4233 6469 4236
rect 6503 4233 6515 4267
rect 8938 4264 8944 4276
rect 8899 4236 8944 4264
rect 6457 4227 6515 4233
rect 8938 4224 8944 4236
rect 8996 4264 9002 4276
rect 9582 4264 9588 4276
rect 8996 4236 9588 4264
rect 8996 4224 9002 4236
rect 9582 4224 9588 4236
rect 9640 4224 9646 4276
rect 12710 4224 12716 4276
rect 12768 4264 12774 4276
rect 12894 4264 12900 4276
rect 12768 4236 12900 4264
rect 12768 4224 12774 4236
rect 12894 4224 12900 4236
rect 12952 4224 12958 4276
rect 14458 4264 14464 4276
rect 14419 4236 14464 4264
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 4338 4196 4344 4208
rect 4299 4168 4344 4196
rect 4338 4156 4344 4168
rect 4396 4156 4402 4208
rect 6178 4156 6184 4208
rect 6236 4196 6242 4208
rect 9306 4196 9312 4208
rect 6236 4168 6592 4196
rect 6236 4156 6242 4168
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 2188 4100 2233 4128
rect 2188 4088 2194 4100
rect 2406 4088 2412 4140
rect 2464 4128 2470 4140
rect 3237 4131 3295 4137
rect 2464 4100 2509 4128
rect 2464 4088 2470 4100
rect 3237 4097 3249 4131
rect 3283 4097 3295 4131
rect 3970 4128 3976 4140
rect 3931 4100 3976 4128
rect 3237 4091 3295 4097
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 2958 4060 2964 4072
rect 2363 4032 2964 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3252 3992 3280 4091
rect 3970 4088 3976 4100
rect 4028 4128 4034 4140
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 4028 4100 4261 4128
rect 4028 4088 4034 4100
rect 4249 4097 4261 4100
rect 4295 4097 4307 4131
rect 4249 4091 4307 4097
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4060 3939 4063
rect 4356 4060 4384 4156
rect 6564 4137 6592 4168
rect 8864 4168 9312 4196
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 5491 4100 5733 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 5721 4097 5733 4100
rect 5767 4128 5779 4131
rect 6549 4131 6607 4137
rect 5767 4100 6316 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 3927 4032 4384 4060
rect 5353 4063 5411 4069
rect 3927 4029 3939 4032
rect 3881 4023 3939 4029
rect 5353 4029 5365 4063
rect 5399 4060 5411 4063
rect 5813 4063 5871 4069
rect 5813 4060 5825 4063
rect 5399 4032 5825 4060
rect 5399 4029 5411 4032
rect 5353 4023 5411 4029
rect 5813 4029 5825 4032
rect 5859 4029 5871 4063
rect 6288 4060 6316 4100
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 7006 4128 7012 4140
rect 6967 4100 7012 4128
rect 6549 4091 6607 4097
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7098 4088 7104 4140
rect 7156 4128 7162 4140
rect 7285 4131 7343 4137
rect 7285 4128 7297 4131
rect 7156 4100 7297 4128
rect 7156 4088 7162 4100
rect 7285 4097 7297 4100
rect 7331 4097 7343 4131
rect 7285 4091 7343 4097
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 8202 4128 8208 4140
rect 8163 4100 8208 4128
rect 7377 4091 7435 4097
rect 7116 4060 7144 4088
rect 6288 4032 7144 4060
rect 7392 4060 7420 4091
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4128 8447 4131
rect 8662 4128 8668 4140
rect 8435 4100 8668 4128
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 8864 4137 8892 4168
rect 9306 4156 9312 4168
rect 9364 4156 9370 4208
rect 11885 4199 11943 4205
rect 11885 4165 11897 4199
rect 11931 4196 11943 4199
rect 12802 4196 12808 4208
rect 11931 4168 12808 4196
rect 11931 4165 11943 4168
rect 11885 4159 11943 4165
rect 12802 4156 12808 4168
rect 12860 4156 12866 4208
rect 12986 4156 12992 4208
rect 13044 4196 13050 4208
rect 13081 4199 13139 4205
rect 13081 4196 13093 4199
rect 13044 4168 13093 4196
rect 13044 4156 13050 4168
rect 13081 4165 13093 4168
rect 13127 4165 13139 4199
rect 13081 4159 13139 4165
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4128 9091 4131
rect 9122 4128 9128 4140
rect 9079 4100 9128 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 9272 4100 9505 4128
rect 9272 4088 9278 4100
rect 9493 4097 9505 4100
rect 9539 4097 9551 4131
rect 10134 4128 10140 4140
rect 10095 4100 10140 4128
rect 9493 4091 9551 4097
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4128 11023 4131
rect 11698 4128 11704 4140
rect 11011 4100 11704 4128
rect 11011 4097 11023 4100
rect 10965 4091 11023 4097
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4128 11851 4131
rect 11974 4128 11980 4140
rect 11839 4100 11980 4128
rect 11839 4097 11851 4100
rect 11793 4091 11851 4097
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 12069 4131 12127 4137
rect 12069 4097 12081 4131
rect 12115 4097 12127 4131
rect 12069 4091 12127 4097
rect 10873 4063 10931 4069
rect 7392 4032 9536 4060
rect 5813 4023 5871 4029
rect 5718 3992 5724 4004
rect 3252 3964 5724 3992
rect 5718 3952 5724 3964
rect 5776 3952 5782 4004
rect 5828 3992 5856 4023
rect 7101 3995 7159 4001
rect 5828 3964 6592 3992
rect 1857 3927 1915 3933
rect 1857 3893 1869 3927
rect 1903 3924 1915 3927
rect 2958 3924 2964 3936
rect 1903 3896 2964 3924
rect 1903 3893 1915 3896
rect 1857 3887 1915 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 3145 3927 3203 3933
rect 3145 3893 3157 3927
rect 3191 3924 3203 3927
rect 5074 3924 5080 3936
rect 3191 3896 5080 3924
rect 3191 3893 3203 3896
rect 3145 3887 3203 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 6564 3924 6592 3964
rect 7101 3961 7113 3995
rect 7147 3992 7159 3995
rect 7282 3992 7288 4004
rect 7147 3964 7288 3992
rect 7147 3961 7159 3964
rect 7101 3955 7159 3961
rect 7282 3952 7288 3964
rect 7340 3952 7346 4004
rect 7392 3924 7420 4032
rect 8389 3995 8447 4001
rect 8389 3961 8401 3995
rect 8435 3992 8447 3995
rect 9398 3992 9404 4004
rect 8435 3964 9404 3992
rect 8435 3961 8447 3964
rect 8389 3955 8447 3961
rect 9398 3952 9404 3964
rect 9456 3952 9462 4004
rect 9508 3992 9536 4032
rect 10873 4029 10885 4063
rect 10919 4060 10931 4063
rect 11882 4060 11888 4072
rect 10919 4032 11888 4060
rect 10919 4029 10931 4032
rect 10873 4023 10931 4029
rect 11882 4020 11888 4032
rect 11940 4060 11946 4072
rect 12084 4060 12112 4091
rect 12618 4088 12624 4140
rect 12676 4128 12682 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12676 4100 12909 4128
rect 12676 4088 12682 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 13354 4088 13360 4140
rect 13412 4128 13418 4140
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13412 4100 13829 4128
rect 13412 4088 13418 4100
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 14182 4128 14188 4140
rect 14143 4100 14188 4128
rect 13817 4091 13875 4097
rect 14182 4088 14188 4100
rect 14240 4088 14246 4140
rect 14274 4088 14280 4140
rect 14332 4128 14338 4140
rect 14642 4128 14648 4140
rect 14332 4100 14648 4128
rect 14332 4088 14338 4100
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 11940 4032 12112 4060
rect 13265 4063 13323 4069
rect 11940 4020 11946 4032
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13538 4060 13544 4072
rect 13311 4032 13544 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 13538 4020 13544 4032
rect 13596 4060 13602 4072
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 13596 4032 14013 4060
rect 13596 4020 13602 4032
rect 14001 4029 14013 4032
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 14093 4063 14151 4069
rect 14093 4029 14105 4063
rect 14139 4029 14151 4063
rect 14093 4023 14151 4029
rect 11517 3995 11575 4001
rect 11517 3992 11529 3995
rect 9508 3964 11529 3992
rect 11517 3961 11529 3964
rect 11563 3961 11575 3995
rect 11517 3955 11575 3961
rect 11974 3952 11980 4004
rect 12032 3992 12038 4004
rect 13446 3992 13452 4004
rect 12032 3964 13452 3992
rect 12032 3952 12038 3964
rect 13446 3952 13452 3964
rect 13504 3952 13510 4004
rect 13906 3952 13912 4004
rect 13964 3992 13970 4004
rect 14108 3992 14136 4023
rect 13964 3964 14136 3992
rect 13964 3952 13970 3964
rect 6564 3896 7420 3924
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7561 3927 7619 3933
rect 7561 3924 7573 3927
rect 7524 3896 7573 3924
rect 7524 3884 7530 3896
rect 7561 3893 7573 3896
rect 7607 3893 7619 3927
rect 9582 3924 9588 3936
rect 9543 3896 9588 3924
rect 7561 3887 7619 3893
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 10229 3927 10287 3933
rect 10229 3893 10241 3927
rect 10275 3924 10287 3927
rect 11238 3924 11244 3936
rect 10275 3896 11244 3924
rect 10275 3893 10287 3896
rect 10229 3887 10287 3893
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 1104 3834 15732 3856
rect 1104 3782 3420 3834
rect 3472 3782 3484 3834
rect 3536 3782 3548 3834
rect 3600 3782 3612 3834
rect 3664 3782 8296 3834
rect 8348 3782 8360 3834
rect 8412 3782 8424 3834
rect 8476 3782 8488 3834
rect 8540 3782 13172 3834
rect 13224 3782 13236 3834
rect 13288 3782 13300 3834
rect 13352 3782 13364 3834
rect 13416 3782 15732 3834
rect 1104 3760 15732 3782
rect 12618 3720 12624 3732
rect 2746 3692 12624 3720
rect 2133 3655 2191 3661
rect 2133 3621 2145 3655
rect 2179 3652 2191 3655
rect 2746 3652 2774 3692
rect 12618 3680 12624 3692
rect 12676 3680 12682 3732
rect 14090 3720 14096 3732
rect 14051 3692 14096 3720
rect 14090 3680 14096 3692
rect 14148 3680 14154 3732
rect 5074 3652 5080 3664
rect 2179 3624 2774 3652
rect 5035 3624 5080 3652
rect 2179 3621 2191 3624
rect 2133 3615 2191 3621
rect 5074 3612 5080 3624
rect 5132 3612 5138 3664
rect 6365 3655 6423 3661
rect 6365 3621 6377 3655
rect 6411 3652 6423 3655
rect 6454 3652 6460 3664
rect 6411 3624 6460 3652
rect 6411 3621 6423 3624
rect 6365 3615 6423 3621
rect 6454 3612 6460 3624
rect 6512 3612 6518 3664
rect 6840 3624 7788 3652
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 2409 3587 2467 3593
rect 2409 3584 2421 3587
rect 1903 3556 2421 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 2409 3553 2421 3556
rect 2455 3584 2467 3587
rect 2774 3584 2780 3596
rect 2455 3556 2780 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 4617 3587 4675 3593
rect 4617 3553 4629 3587
rect 4663 3584 4675 3587
rect 4982 3584 4988 3596
rect 4663 3556 4988 3584
rect 4663 3553 4675 3556
rect 4617 3547 4675 3553
rect 4982 3544 4988 3556
rect 5040 3584 5046 3596
rect 6840 3584 6868 3624
rect 5040 3556 6868 3584
rect 5040 3544 5046 3556
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 6972 3556 7113 3584
rect 6972 3544 6978 3556
rect 7101 3553 7113 3556
rect 7147 3584 7159 3587
rect 7650 3584 7656 3596
rect 7147 3556 7656 3584
rect 7147 3553 7159 3556
rect 7101 3547 7159 3553
rect 7650 3544 7656 3556
rect 7708 3544 7714 3596
rect 7760 3584 7788 3624
rect 8662 3612 8668 3664
rect 8720 3652 8726 3664
rect 9677 3655 9735 3661
rect 9677 3652 9689 3655
rect 8720 3624 9689 3652
rect 8720 3612 8726 3624
rect 9677 3621 9689 3624
rect 9723 3652 9735 3655
rect 12710 3652 12716 3664
rect 9723 3624 12716 3652
rect 9723 3621 9735 3624
rect 9677 3615 9735 3621
rect 12710 3612 12716 3624
rect 12768 3652 12774 3664
rect 14369 3655 14427 3661
rect 14369 3652 14381 3655
rect 12768 3624 14381 3652
rect 12768 3612 12774 3624
rect 14369 3621 14381 3624
rect 14415 3621 14427 3655
rect 14369 3615 14427 3621
rect 9582 3584 9588 3596
rect 7760 3556 9168 3584
rect 9543 3556 9588 3584
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 3234 3516 3240 3528
rect 2087 3488 2360 3516
rect 3147 3488 3240 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 2332 3389 2360 3488
rect 3234 3476 3240 3488
rect 3292 3516 3298 3528
rect 3694 3516 3700 3528
rect 3292 3488 3700 3516
rect 3292 3476 3298 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 3970 3516 3976 3528
rect 3931 3488 3976 3516
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 4798 3516 4804 3528
rect 4759 3488 4804 3516
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5350 3516 5356 3528
rect 5215 3488 5356 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 3602 3408 3608 3460
rect 3660 3448 3666 3460
rect 3881 3451 3939 3457
rect 3881 3448 3893 3451
rect 3660 3420 3893 3448
rect 3660 3408 3666 3420
rect 3881 3417 3893 3420
rect 3927 3417 3939 3451
rect 3881 3411 3939 3417
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 4908 3448 4936 3479
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3516 6239 3519
rect 6362 3516 6368 3528
rect 6227 3488 6368 3516
rect 6227 3485 6239 3488
rect 6181 3479 6239 3485
rect 6362 3476 6368 3488
rect 6420 3476 6426 3528
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6932 3516 6960 3544
rect 6512 3488 6960 3516
rect 6512 3476 6518 3488
rect 7006 3476 7012 3528
rect 7064 3516 7070 3528
rect 7190 3516 7196 3528
rect 7064 3488 7109 3516
rect 7151 3488 7196 3516
rect 7064 3476 7070 3488
rect 7190 3476 7196 3488
rect 7248 3476 7254 3528
rect 7282 3476 7288 3528
rect 7340 3516 7346 3528
rect 7466 3516 7472 3528
rect 7340 3488 7385 3516
rect 7427 3488 7472 3516
rect 7340 3476 7346 3488
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 7935 3519 7993 3525
rect 7935 3518 7947 3519
rect 7852 3490 7947 3518
rect 4212 3420 4936 3448
rect 5368 3448 5396 3476
rect 5368 3420 6868 3448
rect 4212 3408 4218 3420
rect 2317 3383 2375 3389
rect 2317 3349 2329 3383
rect 2363 3380 2375 3383
rect 2958 3380 2964 3392
rect 2363 3352 2964 3380
rect 2363 3349 2375 3352
rect 2317 3343 2375 3349
rect 2958 3340 2964 3352
rect 3016 3340 3022 3392
rect 3145 3383 3203 3389
rect 3145 3349 3157 3383
rect 3191 3380 3203 3383
rect 3786 3380 3792 3392
rect 3191 3352 3792 3380
rect 3191 3349 3203 3352
rect 3145 3343 3203 3349
rect 3786 3340 3792 3352
rect 3844 3340 3850 3392
rect 6840 3389 6868 3420
rect 7650 3408 7656 3460
rect 7708 3448 7714 3460
rect 7852 3448 7880 3490
rect 7935 3485 7947 3490
rect 7981 3485 7993 3519
rect 7935 3479 7993 3485
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 8754 3516 8760 3528
rect 8168 3488 8760 3516
rect 8168 3476 8174 3488
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 7708 3420 7880 3448
rect 7708 3408 7714 3420
rect 6825 3383 6883 3389
rect 6825 3349 6837 3383
rect 6871 3349 6883 3383
rect 6825 3343 6883 3349
rect 7098 3340 7104 3392
rect 7156 3380 7162 3392
rect 7834 3380 7840 3392
rect 7156 3352 7840 3380
rect 7156 3340 7162 3352
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 8018 3380 8024 3392
rect 7979 3352 8024 3380
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 9140 3380 9168 3556
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 9858 3544 9864 3596
rect 9916 3544 9922 3596
rect 9953 3587 10011 3593
rect 9953 3553 9965 3587
rect 9999 3584 10011 3587
rect 11977 3587 12035 3593
rect 9999 3556 11928 3584
rect 9999 3553 10011 3556
rect 9953 3547 10011 3553
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 9493 3519 9551 3525
rect 9493 3485 9505 3519
rect 9539 3516 9551 3519
rect 9674 3516 9680 3528
rect 9539 3488 9680 3516
rect 9539 3485 9551 3488
rect 9493 3479 9551 3485
rect 9324 3448 9352 3479
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3516 9827 3519
rect 9876 3516 9904 3544
rect 11900 3528 11928 3556
rect 11977 3553 11989 3587
rect 12023 3584 12035 3587
rect 12894 3584 12900 3596
rect 12023 3556 12900 3584
rect 12023 3553 12035 3556
rect 11977 3547 12035 3553
rect 12894 3544 12900 3556
rect 12952 3544 12958 3596
rect 14458 3584 14464 3596
rect 14419 3556 14464 3584
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 14553 3587 14611 3593
rect 14553 3553 14565 3587
rect 14599 3584 14611 3587
rect 14599 3556 14872 3584
rect 14599 3553 14611 3556
rect 14553 3547 14611 3553
rect 9815 3488 9904 3516
rect 9815 3485 9827 3488
rect 9769 3479 9827 3485
rect 10134 3476 10140 3528
rect 10192 3516 10198 3528
rect 10873 3519 10931 3525
rect 10873 3516 10885 3519
rect 10192 3488 10885 3516
rect 10192 3476 10198 3488
rect 10873 3485 10885 3488
rect 10919 3485 10931 3519
rect 11054 3516 11060 3528
rect 11015 3488 11060 3516
rect 10873 3479 10931 3485
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 11238 3516 11244 3528
rect 11199 3488 11244 3516
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 11882 3516 11888 3528
rect 11795 3488 11888 3516
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 12161 3519 12219 3525
rect 12161 3485 12173 3519
rect 12207 3485 12219 3519
rect 12161 3479 12219 3485
rect 9858 3448 9864 3460
rect 9324 3420 9864 3448
rect 9858 3408 9864 3420
rect 9916 3408 9922 3460
rect 11146 3448 11152 3460
rect 11107 3420 11152 3448
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 12176 3448 12204 3479
rect 12250 3476 12256 3528
rect 12308 3516 12314 3528
rect 13357 3519 13415 3525
rect 12308 3488 12353 3516
rect 12308 3476 12314 3488
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 13998 3516 14004 3528
rect 13403 3488 14004 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 14274 3516 14280 3528
rect 14235 3488 14280 3516
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 14642 3476 14648 3528
rect 14700 3516 14706 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14700 3488 14749 3516
rect 14700 3476 14706 3488
rect 14737 3485 14749 3488
rect 14783 3485 14795 3519
rect 14737 3479 14795 3485
rect 13538 3448 13544 3460
rect 11256 3420 12204 3448
rect 13499 3420 13544 3448
rect 11256 3380 11284 3420
rect 13538 3408 13544 3420
rect 13596 3408 13602 3460
rect 14844 3448 14872 3556
rect 13648 3420 14872 3448
rect 13648 3392 13676 3420
rect 9140 3352 11284 3380
rect 11425 3383 11483 3389
rect 11425 3349 11437 3383
rect 11471 3380 11483 3383
rect 11790 3380 11796 3392
rect 11471 3352 11796 3380
rect 11471 3349 11483 3352
rect 11425 3343 11483 3349
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 12437 3383 12495 3389
rect 12437 3349 12449 3383
rect 12483 3380 12495 3383
rect 13630 3380 13636 3392
rect 12483 3352 13636 3380
rect 12483 3349 12495 3352
rect 12437 3343 12495 3349
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 1104 3290 15732 3312
rect 1104 3238 5858 3290
rect 5910 3238 5922 3290
rect 5974 3238 5986 3290
rect 6038 3238 6050 3290
rect 6102 3238 10734 3290
rect 10786 3238 10798 3290
rect 10850 3238 10862 3290
rect 10914 3238 10926 3290
rect 10978 3238 15732 3290
rect 1104 3216 15732 3238
rect 7098 3176 7104 3188
rect 2746 3148 7104 3176
rect 1394 2972 1400 2984
rect 1355 2944 1400 2972
rect 1394 2932 1400 2944
rect 1452 2932 1458 2984
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 2746 2972 2774 3148
rect 7098 3136 7104 3148
rect 7156 3136 7162 3188
rect 7282 3136 7288 3188
rect 7340 3176 7346 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7340 3148 7757 3176
rect 7340 3136 7346 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 8573 3179 8631 3185
rect 8573 3145 8585 3179
rect 8619 3176 8631 3179
rect 8662 3176 8668 3188
rect 8619 3148 8668 3176
rect 8619 3145 8631 3148
rect 8573 3139 8631 3145
rect 3786 3108 3792 3120
rect 3747 3080 3792 3108
rect 3786 3068 3792 3080
rect 3844 3068 3850 3120
rect 5626 3108 5632 3120
rect 5587 3080 5632 3108
rect 5626 3068 5632 3080
rect 5684 3068 5690 3120
rect 7650 3108 7656 3120
rect 5828 3080 7656 3108
rect 2866 3040 2872 3052
rect 2827 3012 2872 3040
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 3142 3000 3148 3052
rect 3200 3040 3206 3052
rect 3602 3040 3608 3052
rect 3200 3012 3608 3040
rect 3200 3000 3206 3012
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 3970 3040 3976 3052
rect 3752 3012 3797 3040
rect 3883 3012 3976 3040
rect 3752 3000 3758 3012
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 4614 3040 4620 3052
rect 4575 3012 4620 3040
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 5074 3000 5080 3052
rect 5132 3040 5138 3052
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 5132 3012 5457 3040
rect 5132 3000 5138 3012
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 5534 3000 5540 3052
rect 5592 3040 5598 3052
rect 5592 3012 5637 3040
rect 5592 3000 5598 3012
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 5828 3049 5856 3080
rect 7650 3068 7656 3080
rect 7708 3068 7714 3120
rect 7760 3108 7788 3139
rect 8662 3136 8668 3148
rect 8720 3136 8726 3188
rect 9214 3176 9220 3188
rect 9175 3148 9220 3176
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9401 3179 9459 3185
rect 9401 3145 9413 3179
rect 9447 3176 9459 3179
rect 9766 3176 9772 3188
rect 9447 3148 9772 3176
rect 9447 3145 9459 3148
rect 9401 3139 9459 3145
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 10321 3179 10379 3185
rect 10321 3145 10333 3179
rect 10367 3145 10379 3179
rect 10321 3139 10379 3145
rect 10336 3108 10364 3139
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 11514 3176 11520 3188
rect 11204 3148 11520 3176
rect 11204 3136 11210 3148
rect 11514 3136 11520 3148
rect 11572 3176 11578 3188
rect 11609 3179 11667 3185
rect 11609 3176 11621 3179
rect 11572 3148 11621 3176
rect 11572 3136 11578 3148
rect 11609 3145 11621 3148
rect 11655 3145 11667 3179
rect 11609 3139 11667 3145
rect 7760 3080 10364 3108
rect 10873 3111 10931 3117
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 5776 3012 5825 3040
rect 5776 3000 5782 3012
rect 5813 3009 5825 3012
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3040 6791 3043
rect 7285 3043 7343 3049
rect 6779 3012 7236 3040
rect 6779 3009 6791 3012
rect 6733 3003 6791 3009
rect 1719 2944 2774 2972
rect 3988 2972 4016 3000
rect 6822 2972 6828 2984
rect 3988 2944 6828 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 1854 2864 1860 2916
rect 1912 2904 1918 2916
rect 2685 2907 2743 2913
rect 2685 2904 2697 2907
rect 1912 2876 2697 2904
rect 1912 2864 1918 2876
rect 2685 2873 2697 2876
rect 2731 2873 2743 2907
rect 2685 2867 2743 2873
rect 3786 2864 3792 2916
rect 3844 2904 3850 2916
rect 4433 2907 4491 2913
rect 4433 2904 4445 2907
rect 3844 2876 4445 2904
rect 3844 2864 3850 2876
rect 4433 2873 4445 2876
rect 4479 2873 4491 2907
rect 4433 2867 4491 2873
rect 5166 2864 5172 2916
rect 5224 2904 5230 2916
rect 5224 2876 5396 2904
rect 5224 2864 5230 2876
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3421 2839 3479 2845
rect 3421 2836 3433 2839
rect 2832 2808 3433 2836
rect 2832 2796 2838 2808
rect 3421 2805 3433 2808
rect 3467 2805 3479 2839
rect 3421 2799 3479 2805
rect 4338 2796 4344 2848
rect 4396 2836 4402 2848
rect 4798 2836 4804 2848
rect 4396 2808 4804 2836
rect 4396 2796 4402 2808
rect 4798 2796 4804 2808
rect 4856 2836 4862 2848
rect 5261 2839 5319 2845
rect 5261 2836 5273 2839
rect 4856 2808 5273 2836
rect 4856 2796 4862 2808
rect 5261 2805 5273 2808
rect 5307 2805 5319 2839
rect 5368 2836 5396 2876
rect 5534 2864 5540 2916
rect 5592 2904 5598 2916
rect 6549 2907 6607 2913
rect 6549 2904 6561 2907
rect 5592 2876 6561 2904
rect 5592 2864 5598 2876
rect 6549 2873 6561 2876
rect 6595 2873 6607 2907
rect 7098 2904 7104 2916
rect 6549 2867 6607 2873
rect 6656 2876 7104 2904
rect 6656 2836 6684 2876
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 7208 2904 7236 3012
rect 7285 3009 7297 3043
rect 7331 3040 7343 3043
rect 7466 3040 7472 3052
rect 7331 3012 7472 3040
rect 7331 3009 7343 3012
rect 7285 3003 7343 3009
rect 7466 3000 7472 3012
rect 7524 3040 7530 3052
rect 7748 3043 7806 3049
rect 7748 3040 7760 3043
rect 7524 3012 7760 3040
rect 7524 3000 7530 3012
rect 7748 3009 7760 3012
rect 7794 3009 7806 3043
rect 7748 3003 7806 3009
rect 7377 2975 7435 2981
rect 7377 2941 7389 2975
rect 7423 2972 7435 2975
rect 7852 2972 7880 3080
rect 10873 3077 10885 3111
rect 10919 3108 10931 3111
rect 11790 3108 11796 3120
rect 10919 3080 11796 3108
rect 10919 3077 10931 3080
rect 10873 3071 10931 3077
rect 8665 3043 8723 3049
rect 8665 3009 8677 3043
rect 8711 3040 8723 3043
rect 9030 3040 9036 3052
rect 8711 3012 9036 3040
rect 8711 3009 8723 3012
rect 8665 3003 8723 3009
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 9398 3043 9456 3049
rect 9398 3009 9410 3043
rect 9444 3040 9456 3043
rect 10597 3043 10655 3049
rect 9444 3012 9904 3040
rect 9444 3009 9456 3012
rect 9398 3003 9456 3009
rect 9876 2984 9904 3012
rect 10597 3009 10609 3043
rect 10643 3040 10655 3043
rect 10888 3040 10916 3071
rect 11790 3068 11796 3080
rect 11848 3068 11854 3120
rect 13648 3080 14504 3108
rect 13648 3052 13676 3080
rect 10643 3012 10916 3040
rect 10643 3009 10655 3012
rect 10597 3003 10655 3009
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11112 3012 11529 3040
rect 11112 3000 11118 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 11882 3000 11888 3052
rect 11940 3040 11946 3052
rect 12161 3043 12219 3049
rect 12161 3040 12173 3043
rect 11940 3012 12173 3040
rect 11940 3000 11946 3012
rect 12161 3009 12173 3012
rect 12207 3009 12219 3043
rect 12161 3003 12219 3009
rect 12345 3043 12403 3049
rect 12345 3009 12357 3043
rect 12391 3040 12403 3043
rect 12894 3040 12900 3052
rect 12391 3012 12900 3040
rect 12391 3009 12403 3012
rect 12345 3003 12403 3009
rect 7423 2944 7880 2972
rect 7423 2941 7435 2944
rect 7377 2935 7435 2941
rect 7926 2932 7932 2984
rect 7984 2972 7990 2984
rect 9858 2972 9864 2984
rect 7984 2944 9076 2972
rect 9819 2944 9864 2972
rect 7984 2932 7990 2944
rect 8938 2904 8944 2916
rect 7208 2876 8944 2904
rect 8938 2864 8944 2876
rect 8996 2864 9002 2916
rect 9048 2904 9076 2944
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 10965 2975 11023 2981
rect 10965 2972 10977 2975
rect 10551 2944 10977 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 10965 2941 10977 2944
rect 11011 2972 11023 2975
rect 11974 2972 11980 2984
rect 11011 2944 11980 2972
rect 11011 2941 11023 2944
rect 10965 2935 11023 2941
rect 11974 2932 11980 2944
rect 12032 2932 12038 2984
rect 12176 2972 12204 3003
rect 12894 3000 12900 3012
rect 12952 3040 12958 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12952 3012 13001 3040
rect 12952 3000 12958 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 13630 3040 13636 3052
rect 13591 3012 13636 3040
rect 12989 3003 13047 3009
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 14476 3049 14504 3080
rect 14001 3043 14059 3049
rect 14001 3009 14013 3043
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 14461 3043 14519 3049
rect 14461 3009 14473 3043
rect 14507 3009 14519 3043
rect 14461 3003 14519 3009
rect 13081 2975 13139 2981
rect 13081 2972 13093 2975
rect 12176 2944 13093 2972
rect 13081 2941 13093 2944
rect 13127 2941 13139 2975
rect 14016 2972 14044 3003
rect 14642 2972 14648 2984
rect 14016 2944 14648 2972
rect 13081 2935 13139 2941
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 9950 2904 9956 2916
rect 9048 2876 9956 2904
rect 9950 2864 9956 2876
rect 10008 2864 10014 2916
rect 11146 2864 11152 2916
rect 11204 2904 11210 2916
rect 12250 2904 12256 2916
rect 11204 2876 12256 2904
rect 11204 2864 11210 2876
rect 12250 2864 12256 2876
rect 12308 2904 12314 2916
rect 12437 2907 12495 2913
rect 12437 2904 12449 2907
rect 12308 2876 12449 2904
rect 12308 2864 12314 2876
rect 12437 2873 12449 2876
rect 12483 2873 12495 2907
rect 12437 2867 12495 2873
rect 14185 2907 14243 2913
rect 14185 2873 14197 2907
rect 14231 2873 14243 2907
rect 14185 2867 14243 2873
rect 5368 2808 6684 2836
rect 5261 2799 5319 2805
rect 6730 2796 6736 2848
rect 6788 2836 6794 2848
rect 7374 2836 7380 2848
rect 6788 2808 7380 2836
rect 6788 2796 6794 2808
rect 7374 2796 7380 2808
rect 7432 2796 7438 2848
rect 7926 2836 7932 2848
rect 7887 2808 7932 2836
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 9122 2796 9128 2848
rect 9180 2836 9186 2848
rect 9490 2836 9496 2848
rect 9180 2808 9496 2836
rect 9180 2796 9186 2808
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 9766 2836 9772 2848
rect 9679 2808 9772 2836
rect 9766 2796 9772 2808
rect 9824 2836 9830 2848
rect 12066 2836 12072 2848
rect 9824 2808 12072 2836
rect 9824 2796 9830 2808
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 12158 2796 12164 2848
rect 12216 2836 12222 2848
rect 14200 2836 14228 2867
rect 12216 2808 14228 2836
rect 12216 2796 12222 2808
rect 1104 2746 15732 2768
rect 1104 2694 3420 2746
rect 3472 2694 3484 2746
rect 3536 2694 3548 2746
rect 3600 2694 3612 2746
rect 3664 2694 8296 2746
rect 8348 2694 8360 2746
rect 8412 2694 8424 2746
rect 8476 2694 8488 2746
rect 8540 2694 13172 2746
rect 13224 2694 13236 2746
rect 13288 2694 13300 2746
rect 13352 2694 13364 2746
rect 13416 2694 15732 2746
rect 1104 2672 15732 2694
rect 3142 2632 3148 2644
rect 3103 2604 3148 2632
rect 3142 2592 3148 2604
rect 3200 2592 3206 2644
rect 4614 2592 4620 2644
rect 4672 2632 4678 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 4672 2604 5089 2632
rect 4672 2592 4678 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 5077 2595 5135 2601
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 8021 2635 8079 2641
rect 8021 2632 8033 2635
rect 7248 2604 8033 2632
rect 7248 2592 7254 2604
rect 8021 2601 8033 2604
rect 8067 2601 8079 2635
rect 11146 2632 11152 2644
rect 8021 2595 8079 2601
rect 9232 2604 11152 2632
rect 2866 2524 2872 2576
rect 2924 2564 2930 2576
rect 4065 2567 4123 2573
rect 4065 2564 4077 2567
rect 2924 2536 4077 2564
rect 2924 2524 2930 2536
rect 4065 2533 4077 2536
rect 4111 2533 4123 2567
rect 4065 2527 4123 2533
rect 6914 2524 6920 2576
rect 6972 2564 6978 2576
rect 7101 2567 7159 2573
rect 7101 2564 7113 2567
rect 6972 2536 7113 2564
rect 6972 2524 6978 2536
rect 7101 2533 7113 2536
rect 7147 2564 7159 2567
rect 9030 2564 9036 2576
rect 7147 2536 9036 2564
rect 7147 2533 7159 2536
rect 7101 2527 7159 2533
rect 9030 2524 9036 2536
rect 9088 2524 9094 2576
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 3050 2496 3056 2508
rect 1719 2468 3056 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 3050 2456 3056 2468
rect 3108 2456 3114 2508
rect 3789 2499 3847 2505
rect 3789 2465 3801 2499
rect 3835 2496 3847 2499
rect 4338 2496 4344 2508
rect 3835 2468 4344 2496
rect 3835 2465 3847 2468
rect 3789 2459 3847 2465
rect 4338 2456 4344 2468
rect 4396 2456 4402 2508
rect 4801 2499 4859 2505
rect 4801 2465 4813 2499
rect 4847 2496 4859 2499
rect 5353 2499 5411 2505
rect 5353 2496 5365 2499
rect 4847 2468 5365 2496
rect 4847 2465 4859 2468
rect 4801 2459 4859 2465
rect 5353 2465 5365 2468
rect 5399 2496 5411 2499
rect 7190 2496 7196 2508
rect 5399 2468 6914 2496
rect 7151 2468 7196 2496
rect 5399 2465 5411 2468
rect 5353 2459 5411 2465
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2832 2400 2881 2428
rect 2832 2388 2838 2400
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 2958 2388 2964 2440
rect 3016 2428 3022 2440
rect 3234 2428 3240 2440
rect 3016 2400 3061 2428
rect 3195 2400 3240 2428
rect 3016 2388 3022 2400
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 4154 2428 4160 2440
rect 3896 2400 4160 2428
rect 3896 2369 3924 2400
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 2685 2363 2743 2369
rect 2685 2329 2697 2363
rect 2731 2360 2743 2363
rect 3881 2363 3939 2369
rect 3881 2360 3893 2363
rect 2731 2332 3893 2360
rect 2731 2329 2743 2332
rect 2685 2323 2743 2329
rect 3881 2329 3893 2332
rect 3927 2329 3939 2363
rect 3881 2323 3939 2329
rect 4893 2363 4951 2369
rect 4893 2329 4905 2363
rect 4939 2360 4951 2363
rect 4982 2360 4988 2372
rect 4939 2332 4988 2360
rect 4939 2329 4951 2332
rect 4893 2323 4951 2329
rect 4982 2320 4988 2332
rect 5040 2360 5046 2372
rect 5184 2360 5212 2391
rect 5040 2332 5212 2360
rect 6886 2360 6914 2468
rect 7190 2456 7196 2468
rect 7248 2456 7254 2508
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 8018 2496 8024 2508
rect 7331 2468 8024 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 8018 2456 8024 2468
rect 8076 2456 8082 2508
rect 9232 2496 9260 2604
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11238 2592 11244 2644
rect 11296 2632 11302 2644
rect 11609 2635 11667 2641
rect 11609 2632 11621 2635
rect 11296 2604 11621 2632
rect 11296 2592 11302 2604
rect 11609 2601 11621 2604
rect 11655 2601 11667 2635
rect 11609 2595 11667 2601
rect 12526 2592 12532 2644
rect 12584 2632 12590 2644
rect 13357 2635 13415 2641
rect 13357 2632 13369 2635
rect 12584 2604 13369 2632
rect 12584 2592 12590 2604
rect 13357 2601 13369 2604
rect 13403 2601 13415 2635
rect 13357 2595 13415 2601
rect 14642 2592 14648 2644
rect 14700 2632 14706 2644
rect 15013 2635 15071 2641
rect 15013 2632 15025 2635
rect 14700 2604 15025 2632
rect 14700 2592 14706 2604
rect 15013 2601 15025 2604
rect 15059 2601 15071 2635
rect 15013 2595 15071 2601
rect 9582 2524 9588 2576
rect 9640 2524 9646 2576
rect 9858 2524 9864 2576
rect 9916 2564 9922 2576
rect 12069 2567 12127 2573
rect 12069 2564 12081 2567
rect 9916 2536 12081 2564
rect 9916 2524 9922 2536
rect 12069 2533 12081 2536
rect 12115 2533 12127 2567
rect 13722 2564 13728 2576
rect 12069 2527 12127 2533
rect 12544 2536 13728 2564
rect 8956 2468 9260 2496
rect 9309 2499 9367 2505
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7469 2431 7527 2437
rect 7064 2400 7109 2428
rect 7064 2388 7070 2400
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7926 2428 7932 2440
rect 7515 2400 7932 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 8956 2360 8984 2468
rect 9309 2465 9321 2499
rect 9355 2496 9367 2499
rect 9600 2496 9628 2524
rect 9355 2468 9628 2496
rect 10873 2499 10931 2505
rect 9355 2465 9367 2468
rect 9309 2459 9367 2465
rect 10873 2465 10885 2499
rect 10919 2496 10931 2499
rect 12544 2496 12572 2536
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 14366 2524 14372 2576
rect 14424 2564 14430 2576
rect 14826 2564 14832 2576
rect 14424 2536 14832 2564
rect 14424 2524 14430 2536
rect 14826 2524 14832 2536
rect 14884 2524 14890 2576
rect 10919 2468 12572 2496
rect 12805 2499 12863 2505
rect 10919 2465 10931 2468
rect 10873 2459 10931 2465
rect 12805 2465 12817 2499
rect 12851 2496 12863 2499
rect 14918 2496 14924 2508
rect 12851 2468 14924 2496
rect 12851 2465 12863 2468
rect 12805 2459 12863 2465
rect 14918 2456 14924 2468
rect 14976 2456 14982 2508
rect 9122 2428 9128 2440
rect 9083 2400 9128 2428
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2397 9275 2431
rect 9398 2428 9404 2440
rect 9359 2400 9404 2428
rect 9217 2391 9275 2397
rect 6886 2332 8984 2360
rect 5040 2320 5046 2332
rect 9030 2320 9036 2372
rect 9088 2360 9094 2372
rect 9232 2360 9260 2391
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2397 11023 2431
rect 11514 2428 11520 2440
rect 11475 2400 11520 2428
rect 10965 2391 11023 2397
rect 9088 2332 9260 2360
rect 9088 2320 9094 2332
rect 9306 2320 9312 2372
rect 9364 2360 9370 2372
rect 9600 2360 9628 2391
rect 10226 2360 10232 2372
rect 9364 2332 9628 2360
rect 10187 2332 10232 2360
rect 9364 2320 9370 2332
rect 10226 2320 10232 2332
rect 10284 2320 10290 2372
rect 10980 2360 11008 2391
rect 11514 2388 11520 2400
rect 11572 2388 11578 2440
rect 11790 2428 11796 2440
rect 11751 2400 11796 2428
rect 11790 2388 11796 2400
rect 11848 2388 11854 2440
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2428 11943 2431
rect 11974 2428 11980 2440
rect 11931 2400 11980 2428
rect 11931 2397 11943 2400
rect 11885 2391 11943 2397
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 12618 2428 12624 2440
rect 12579 2400 12624 2428
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2428 13507 2431
rect 14734 2428 14740 2440
rect 13495 2400 14596 2428
rect 14695 2400 14740 2428
rect 13495 2397 13507 2400
rect 13449 2391 13507 2397
rect 13906 2360 13912 2372
rect 10980 2332 13912 2360
rect 13906 2320 13912 2332
rect 13964 2320 13970 2372
rect 14366 2360 14372 2372
rect 14327 2332 14372 2360
rect 14366 2320 14372 2332
rect 14424 2320 14430 2372
rect 14461 2363 14519 2369
rect 14461 2329 14473 2363
rect 14507 2329 14519 2363
rect 14568 2360 14596 2400
rect 14734 2388 14740 2400
rect 14792 2388 14798 2440
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 14884 2400 14929 2428
rect 14884 2388 14890 2400
rect 16758 2360 16764 2372
rect 14568 2332 16764 2360
rect 14461 2323 14519 2329
rect 6822 2292 6828 2304
rect 6783 2264 6828 2292
rect 6822 2252 6828 2264
rect 6880 2252 6886 2304
rect 7650 2252 7656 2304
rect 7708 2292 7714 2304
rect 8941 2295 8999 2301
rect 8941 2292 8953 2295
rect 7708 2264 8953 2292
rect 7708 2252 7714 2264
rect 8941 2261 8953 2264
rect 8987 2261 8999 2295
rect 8941 2255 8999 2261
rect 9214 2252 9220 2304
rect 9272 2292 9278 2304
rect 10137 2295 10195 2301
rect 10137 2292 10149 2295
rect 9272 2264 10149 2292
rect 9272 2252 9278 2264
rect 10137 2261 10149 2264
rect 10183 2261 10195 2295
rect 14476 2292 14504 2323
rect 16758 2320 16764 2332
rect 16816 2320 16822 2372
rect 14734 2292 14740 2304
rect 14476 2264 14740 2292
rect 10137 2255 10195 2261
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 1104 2202 15732 2224
rect 1104 2150 5858 2202
rect 5910 2150 5922 2202
rect 5974 2150 5986 2202
rect 6038 2150 6050 2202
rect 6102 2150 10734 2202
rect 10786 2150 10798 2202
rect 10850 2150 10862 2202
rect 10914 2150 10926 2202
rect 10978 2150 15732 2202
rect 1104 2128 15732 2150
rect 6638 2048 6644 2100
rect 6696 2088 6702 2100
rect 10226 2088 10232 2100
rect 6696 2060 10232 2088
rect 6696 2048 6702 2060
rect 10226 2048 10232 2060
rect 10284 2048 10290 2100
rect 10594 1912 10600 1964
rect 10652 1952 10658 1964
rect 12894 1952 12900 1964
rect 10652 1924 12900 1952
rect 10652 1912 10658 1924
rect 12894 1912 12900 1924
rect 12952 1912 12958 1964
rect 10502 1096 10508 1148
rect 10560 1136 10566 1148
rect 11054 1136 11060 1148
rect 10560 1108 11060 1136
rect 10560 1096 10566 1108
rect 11054 1096 11060 1108
rect 11112 1096 11118 1148
<< via1 >>
rect 5858 16294 5910 16346
rect 5922 16294 5974 16346
rect 5986 16294 6038 16346
rect 6050 16294 6102 16346
rect 10734 16294 10786 16346
rect 10798 16294 10850 16346
rect 10862 16294 10914 16346
rect 10926 16294 10978 16346
rect 3884 16124 3936 16176
rect 7564 16124 7616 16176
rect 9680 16124 9732 16176
rect 13084 16124 13136 16176
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 2872 16099 2924 16108
rect 2872 16065 2881 16099
rect 2881 16065 2915 16099
rect 2915 16065 2924 16099
rect 2872 16056 2924 16065
rect 2964 16099 3016 16108
rect 2964 16065 2973 16099
rect 2973 16065 3007 16099
rect 3007 16065 3016 16099
rect 3240 16099 3292 16108
rect 2964 16056 3016 16065
rect 3240 16065 3249 16099
rect 3249 16065 3283 16099
rect 3283 16065 3292 16099
rect 3240 16056 3292 16065
rect 4252 16056 4304 16108
rect 5264 16056 5316 16108
rect 5724 16056 5776 16108
rect 9128 16099 9180 16108
rect 6552 15988 6604 16040
rect 6828 15988 6880 16040
rect 9128 16065 9137 16099
rect 9137 16065 9171 16099
rect 9171 16065 9180 16099
rect 9128 16056 9180 16065
rect 9220 16099 9272 16108
rect 9220 16065 9229 16099
rect 9229 16065 9263 16099
rect 9263 16065 9272 16099
rect 9220 16056 9272 16065
rect 9772 16056 9824 16108
rect 10140 16099 10192 16108
rect 10140 16065 10149 16099
rect 10149 16065 10183 16099
rect 10183 16065 10192 16099
rect 10140 16056 10192 16065
rect 11244 16056 11296 16108
rect 16764 16124 16816 16176
rect 14556 16056 14608 16108
rect 14648 16056 14700 16108
rect 15016 16099 15068 16108
rect 15016 16065 15025 16099
rect 15025 16065 15059 16099
rect 15059 16065 15068 16099
rect 15016 16056 15068 16065
rect 12624 15988 12676 16040
rect 4160 15963 4212 15972
rect 4160 15929 4169 15963
rect 4169 15929 4203 15963
rect 4203 15929 4212 15963
rect 4160 15920 4212 15929
rect 13820 15920 13872 15972
rect 2044 15852 2096 15904
rect 3148 15895 3200 15904
rect 3148 15861 3157 15895
rect 3157 15861 3191 15895
rect 3191 15861 3200 15895
rect 3148 15852 3200 15861
rect 5448 15852 5500 15904
rect 9404 15895 9456 15904
rect 9404 15861 9413 15895
rect 9413 15861 9447 15895
rect 9447 15861 9456 15895
rect 9404 15852 9456 15861
rect 11704 15895 11756 15904
rect 11704 15861 11713 15895
rect 11713 15861 11747 15895
rect 11747 15861 11756 15895
rect 11704 15852 11756 15861
rect 12808 15852 12860 15904
rect 14740 15852 14792 15904
rect 3420 15750 3472 15802
rect 3484 15750 3536 15802
rect 3548 15750 3600 15802
rect 3612 15750 3664 15802
rect 8296 15750 8348 15802
rect 8360 15750 8412 15802
rect 8424 15750 8476 15802
rect 8488 15750 8540 15802
rect 13172 15750 13224 15802
rect 13236 15750 13288 15802
rect 13300 15750 13352 15802
rect 13364 15750 13416 15802
rect 9220 15648 9272 15700
rect 14648 15691 14700 15700
rect 14648 15657 14657 15691
rect 14657 15657 14691 15691
rect 14691 15657 14700 15691
rect 14648 15648 14700 15657
rect 2872 15580 2924 15632
rect 1584 15512 1636 15564
rect 2044 15555 2096 15564
rect 2044 15521 2053 15555
rect 2053 15521 2087 15555
rect 2087 15521 2096 15555
rect 2044 15512 2096 15521
rect 5448 15580 5500 15632
rect 12900 15623 12952 15632
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 2964 15444 3016 15496
rect 1860 15351 1912 15360
rect 1860 15317 1869 15351
rect 1869 15317 1903 15351
rect 1903 15317 1912 15351
rect 1860 15308 1912 15317
rect 2872 15308 2924 15360
rect 3424 15308 3476 15360
rect 5632 15376 5684 15428
rect 9404 15512 9456 15564
rect 7380 15444 7432 15496
rect 7932 15487 7984 15496
rect 7932 15453 7941 15487
rect 7941 15453 7975 15487
rect 7975 15453 7984 15487
rect 12900 15589 12909 15623
rect 12909 15589 12943 15623
rect 12943 15589 12952 15623
rect 12900 15580 12952 15589
rect 7932 15444 7984 15453
rect 6184 15419 6236 15428
rect 6184 15385 6193 15419
rect 6193 15385 6227 15419
rect 6227 15385 6236 15419
rect 6184 15376 6236 15385
rect 10416 15444 10468 15496
rect 9772 15376 9824 15428
rect 10324 15376 10376 15428
rect 10508 15419 10560 15428
rect 10508 15385 10517 15419
rect 10517 15385 10551 15419
rect 10551 15385 10560 15419
rect 12072 15444 12124 15496
rect 12256 15419 12308 15428
rect 10508 15376 10560 15385
rect 5356 15308 5408 15360
rect 11796 15351 11848 15360
rect 11796 15317 11805 15351
rect 11805 15317 11839 15351
rect 11839 15317 11848 15351
rect 11796 15308 11848 15317
rect 12256 15385 12265 15419
rect 12265 15385 12299 15419
rect 12299 15385 12308 15419
rect 12992 15444 13044 15496
rect 14188 15444 14240 15496
rect 14280 15444 14332 15496
rect 14464 15419 14516 15428
rect 12256 15376 12308 15385
rect 14004 15308 14056 15360
rect 14464 15385 14473 15419
rect 14473 15385 14507 15419
rect 14507 15385 14516 15419
rect 14464 15376 14516 15385
rect 14924 15308 14976 15360
rect 5858 15206 5910 15258
rect 5922 15206 5974 15258
rect 5986 15206 6038 15258
rect 6050 15206 6102 15258
rect 10734 15206 10786 15258
rect 10798 15206 10850 15258
rect 10862 15206 10914 15258
rect 10926 15206 10978 15258
rect 1952 15104 2004 15156
rect 3424 15147 3476 15156
rect 3424 15113 3433 15147
rect 3433 15113 3467 15147
rect 3467 15113 3476 15147
rect 3424 15104 3476 15113
rect 5356 15147 5408 15156
rect 5356 15113 5365 15147
rect 5365 15113 5399 15147
rect 5399 15113 5408 15147
rect 5356 15104 5408 15113
rect 6184 15104 6236 15156
rect 9220 15104 9272 15156
rect 1860 15036 1912 15088
rect 1584 15011 1636 15020
rect 1584 14977 1593 15011
rect 1593 14977 1627 15011
rect 1627 14977 1636 15011
rect 1584 14968 1636 14977
rect 1676 15011 1728 15020
rect 1676 14977 1685 15011
rect 1685 14977 1719 15011
rect 1719 14977 1728 15011
rect 1676 14968 1728 14977
rect 2044 14968 2096 15020
rect 3148 14968 3200 15020
rect 7932 15036 7984 15088
rect 7380 15011 7432 15020
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7656 15011 7708 15020
rect 7380 14968 7432 14977
rect 7656 14977 7665 15011
rect 7665 14977 7699 15011
rect 7699 14977 7708 15011
rect 7656 14968 7708 14977
rect 10140 15104 10192 15156
rect 12624 15104 12676 15156
rect 14464 15147 14516 15156
rect 14464 15113 14473 15147
rect 14473 15113 14507 15147
rect 14507 15113 14516 15147
rect 14464 15104 14516 15113
rect 3240 14900 3292 14952
rect 4068 14943 4120 14952
rect 4068 14909 4077 14943
rect 4077 14909 4111 14943
rect 4111 14909 4120 14943
rect 4068 14900 4120 14909
rect 5448 14900 5500 14952
rect 9128 14900 9180 14952
rect 20 14832 72 14884
rect 4160 14832 4212 14884
rect 12256 14968 12308 15020
rect 12900 14968 12952 15020
rect 12072 14943 12124 14952
rect 12072 14909 12081 14943
rect 12081 14909 12115 14943
rect 12115 14909 12124 14943
rect 12072 14900 12124 14909
rect 13544 14900 13596 14952
rect 13728 14900 13780 14952
rect 13912 14943 13964 14952
rect 13912 14909 13921 14943
rect 13921 14909 13955 14943
rect 13955 14909 13964 14943
rect 13912 14900 13964 14909
rect 1584 14764 1636 14816
rect 2228 14764 2280 14816
rect 6644 14764 6696 14816
rect 7564 14807 7616 14816
rect 7564 14773 7573 14807
rect 7573 14773 7607 14807
rect 7607 14773 7616 14807
rect 7564 14764 7616 14773
rect 3420 14662 3472 14714
rect 3484 14662 3536 14714
rect 3548 14662 3600 14714
rect 3612 14662 3664 14714
rect 8296 14662 8348 14714
rect 8360 14662 8412 14714
rect 8424 14662 8476 14714
rect 8488 14662 8540 14714
rect 13172 14662 13224 14714
rect 13236 14662 13288 14714
rect 13300 14662 13352 14714
rect 13364 14662 13416 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 4068 14560 4120 14612
rect 7380 14560 7432 14612
rect 7932 14560 7984 14612
rect 10416 14603 10468 14612
rect 10416 14569 10425 14603
rect 10425 14569 10459 14603
rect 10459 14569 10468 14603
rect 10416 14560 10468 14569
rect 12256 14560 12308 14612
rect 13544 14560 13596 14612
rect 5080 14492 5132 14544
rect 2044 14424 2096 14476
rect 7656 14492 7708 14544
rect 2228 14331 2280 14340
rect 2228 14297 2237 14331
rect 2237 14297 2271 14331
rect 2271 14297 2280 14331
rect 2228 14288 2280 14297
rect 4712 14399 4764 14408
rect 4712 14365 4721 14399
rect 4721 14365 4755 14399
rect 4755 14365 4764 14399
rect 4712 14356 4764 14365
rect 4804 14399 4856 14408
rect 4804 14365 4813 14399
rect 4813 14365 4847 14399
rect 4847 14365 4856 14399
rect 4804 14356 4856 14365
rect 5540 14356 5592 14408
rect 12440 14492 12492 14544
rect 13912 14492 13964 14544
rect 2688 14288 2740 14340
rect 7564 14331 7616 14340
rect 7564 14297 7573 14331
rect 7573 14297 7607 14331
rect 7607 14297 7616 14331
rect 7564 14288 7616 14297
rect 9864 14356 9916 14408
rect 4896 14220 4948 14272
rect 7288 14220 7340 14272
rect 8116 14220 8168 14272
rect 9588 14288 9640 14340
rect 12624 14424 12676 14476
rect 13728 14424 13780 14476
rect 11796 14399 11848 14408
rect 11796 14365 11805 14399
rect 11805 14365 11839 14399
rect 11839 14365 11848 14399
rect 11796 14356 11848 14365
rect 12072 14356 12124 14408
rect 12164 14356 12216 14408
rect 12716 14399 12768 14408
rect 12716 14365 12725 14399
rect 12725 14365 12759 14399
rect 12759 14365 12768 14399
rect 12716 14356 12768 14365
rect 12808 14399 12860 14408
rect 12808 14365 12817 14399
rect 12817 14365 12851 14399
rect 12851 14365 12860 14399
rect 14280 14399 14332 14408
rect 12808 14356 12860 14365
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 14464 14356 14516 14408
rect 9404 14220 9456 14272
rect 11060 14331 11112 14340
rect 11060 14297 11069 14331
rect 11069 14297 11103 14331
rect 11103 14297 11112 14331
rect 11060 14288 11112 14297
rect 14740 14288 14792 14340
rect 11152 14220 11204 14272
rect 14372 14220 14424 14272
rect 5858 14118 5910 14170
rect 5922 14118 5974 14170
rect 5986 14118 6038 14170
rect 6050 14118 6102 14170
rect 10734 14118 10786 14170
rect 10798 14118 10850 14170
rect 10862 14118 10914 14170
rect 10926 14118 10978 14170
rect 3148 14059 3200 14068
rect 3148 14025 3157 14059
rect 3157 14025 3191 14059
rect 3191 14025 3200 14059
rect 3148 14016 3200 14025
rect 4804 14059 4856 14068
rect 4804 14025 4813 14059
rect 4813 14025 4847 14059
rect 4847 14025 4856 14059
rect 4804 14016 4856 14025
rect 7564 14016 7616 14068
rect 10324 14059 10376 14068
rect 10324 14025 10333 14059
rect 10333 14025 10367 14059
rect 10367 14025 10376 14059
rect 10324 14016 10376 14025
rect 4896 13948 4948 14000
rect 9312 13948 9364 14000
rect 10416 13948 10468 14000
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 2412 13880 2464 13932
rect 5080 13923 5132 13932
rect 5080 13889 5089 13923
rect 5089 13889 5123 13923
rect 5123 13889 5132 13923
rect 5080 13880 5132 13889
rect 5724 13880 5776 13932
rect 6736 13880 6788 13932
rect 8944 13880 8996 13932
rect 9496 13923 9548 13932
rect 9496 13889 9505 13923
rect 9505 13889 9539 13923
rect 9539 13889 9548 13923
rect 9496 13880 9548 13889
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 3148 13812 3200 13864
rect 5540 13812 5592 13864
rect 5816 13812 5868 13864
rect 8024 13855 8076 13864
rect 8024 13821 8033 13855
rect 8033 13821 8067 13855
rect 8067 13821 8076 13855
rect 8024 13812 8076 13821
rect 11152 13948 11204 14000
rect 11704 13923 11756 13932
rect 11704 13889 11713 13923
rect 11713 13889 11747 13923
rect 11747 13889 11756 13923
rect 11704 13880 11756 13889
rect 12256 13880 12308 13932
rect 12532 13812 12584 13864
rect 12716 13948 12768 14000
rect 13912 14016 13964 14068
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 13544 13812 13596 13864
rect 13820 13880 13872 13932
rect 14832 13923 14884 13932
rect 14832 13889 14841 13923
rect 14841 13889 14875 13923
rect 14875 13889 14884 13923
rect 14832 13880 14884 13889
rect 13912 13812 13964 13864
rect 6184 13744 6236 13796
rect 12808 13744 12860 13796
rect 13636 13744 13688 13796
rect 15016 13855 15068 13864
rect 15016 13821 15025 13855
rect 15025 13821 15059 13855
rect 15059 13821 15068 13855
rect 15016 13812 15068 13821
rect 7104 13719 7156 13728
rect 7104 13685 7113 13719
rect 7113 13685 7147 13719
rect 7147 13685 7156 13719
rect 7104 13676 7156 13685
rect 11060 13676 11112 13728
rect 12624 13676 12676 13728
rect 15108 13676 15160 13728
rect 3420 13574 3472 13626
rect 3484 13574 3536 13626
rect 3548 13574 3600 13626
rect 3612 13574 3664 13626
rect 8296 13574 8348 13626
rect 8360 13574 8412 13626
rect 8424 13574 8476 13626
rect 8488 13574 8540 13626
rect 13172 13574 13224 13626
rect 13236 13574 13288 13626
rect 13300 13574 13352 13626
rect 13364 13574 13416 13626
rect 2688 13515 2740 13524
rect 2688 13481 2697 13515
rect 2697 13481 2731 13515
rect 2731 13481 2740 13515
rect 2688 13472 2740 13481
rect 5632 13472 5684 13524
rect 7196 13515 7248 13524
rect 7196 13481 7205 13515
rect 7205 13481 7239 13515
rect 7239 13481 7248 13515
rect 7196 13472 7248 13481
rect 8024 13472 8076 13524
rect 8944 13515 8996 13524
rect 8944 13481 8953 13515
rect 8953 13481 8987 13515
rect 8987 13481 8996 13515
rect 8944 13472 8996 13481
rect 12532 13515 12584 13524
rect 5816 13404 5868 13456
rect 1676 13336 1728 13388
rect 4804 13336 4856 13388
rect 2412 13311 2464 13320
rect 2412 13277 2421 13311
rect 2421 13277 2455 13311
rect 2455 13277 2464 13311
rect 2412 13268 2464 13277
rect 3148 13268 3200 13320
rect 5356 13311 5408 13320
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 7012 13268 7064 13320
rect 2780 13200 2832 13252
rect 4712 13200 4764 13252
rect 8944 13200 8996 13252
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9220 13268 9272 13277
rect 11888 13336 11940 13388
rect 12532 13481 12541 13515
rect 12541 13481 12575 13515
rect 12575 13481 12584 13515
rect 12532 13472 12584 13481
rect 13544 13472 13596 13524
rect 14740 13515 14792 13524
rect 14740 13481 14749 13515
rect 14749 13481 14783 13515
rect 14783 13481 14792 13515
rect 14740 13472 14792 13481
rect 14188 13404 14240 13456
rect 10232 13268 10284 13320
rect 10600 13268 10652 13320
rect 10876 13268 10928 13320
rect 11336 13311 11388 13320
rect 11336 13277 11345 13311
rect 11345 13277 11379 13311
rect 11379 13277 11388 13311
rect 12164 13336 12216 13388
rect 11336 13268 11388 13277
rect 10048 13200 10100 13252
rect 11888 13243 11940 13252
rect 10324 13175 10376 13184
rect 10324 13141 10333 13175
rect 10333 13141 10367 13175
rect 10367 13141 10376 13175
rect 10324 13132 10376 13141
rect 11888 13209 11897 13243
rect 11897 13209 11931 13243
rect 11931 13209 11940 13243
rect 11888 13200 11940 13209
rect 12164 13200 12216 13252
rect 12440 13268 12492 13320
rect 12900 13268 12952 13320
rect 13636 13268 13688 13320
rect 14096 13268 14148 13320
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 14648 13268 14700 13320
rect 5858 13030 5910 13082
rect 5922 13030 5974 13082
rect 5986 13030 6038 13082
rect 6050 13030 6102 13082
rect 10734 13030 10786 13082
rect 10798 13030 10850 13082
rect 10862 13030 10914 13082
rect 10926 13030 10978 13082
rect 2412 12928 2464 12980
rect 5080 12928 5132 12980
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 3056 12792 3108 12844
rect 8024 12860 8076 12912
rect 10048 12860 10100 12912
rect 1676 12724 1728 12733
rect 2780 12724 2832 12776
rect 5724 12792 5776 12844
rect 6184 12792 6236 12844
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 7104 12792 7156 12844
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 9772 12792 9824 12844
rect 9956 12835 10008 12844
rect 9956 12801 9965 12835
rect 9965 12801 9999 12835
rect 9999 12801 10008 12835
rect 9956 12792 10008 12801
rect 10508 12860 10560 12912
rect 14464 12928 14516 12980
rect 4436 12724 4488 12776
rect 4344 12656 4396 12708
rect 7012 12724 7064 12776
rect 9496 12724 9548 12776
rect 8668 12656 8720 12708
rect 11704 12792 11756 12844
rect 11980 12792 12032 12844
rect 12164 12792 12216 12844
rect 13728 12860 13780 12912
rect 10692 12724 10744 12776
rect 14096 12767 14148 12776
rect 14096 12733 14105 12767
rect 14105 12733 14139 12767
rect 14139 12733 14148 12767
rect 14096 12724 14148 12733
rect 14188 12767 14240 12776
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 14188 12724 14240 12733
rect 4068 12588 4120 12640
rect 6552 12588 6604 12640
rect 8852 12588 8904 12640
rect 10140 12588 10192 12640
rect 11796 12631 11848 12640
rect 11796 12597 11805 12631
rect 11805 12597 11839 12631
rect 11839 12597 11848 12631
rect 11796 12588 11848 12597
rect 12440 12588 12492 12640
rect 3420 12486 3472 12538
rect 3484 12486 3536 12538
rect 3548 12486 3600 12538
rect 3612 12486 3664 12538
rect 8296 12486 8348 12538
rect 8360 12486 8412 12538
rect 8424 12486 8476 12538
rect 8488 12486 8540 12538
rect 13172 12486 13224 12538
rect 13236 12486 13288 12538
rect 13300 12486 13352 12538
rect 13364 12486 13416 12538
rect 2780 12384 2832 12436
rect 5356 12427 5408 12436
rect 5356 12393 5365 12427
rect 5365 12393 5399 12427
rect 5399 12393 5408 12427
rect 5356 12384 5408 12393
rect 7196 12427 7248 12436
rect 7196 12393 7205 12427
rect 7205 12393 7239 12427
rect 7239 12393 7248 12427
rect 7196 12384 7248 12393
rect 7656 12427 7708 12436
rect 7656 12393 7665 12427
rect 7665 12393 7699 12427
rect 7699 12393 7708 12427
rect 7656 12384 7708 12393
rect 8024 12384 8076 12436
rect 8668 12384 8720 12436
rect 9220 12427 9272 12436
rect 9220 12393 9229 12427
rect 9229 12393 9263 12427
rect 9263 12393 9272 12427
rect 9220 12384 9272 12393
rect 8300 12316 8352 12368
rect 4436 12248 4488 12300
rect 7104 12248 7156 12300
rect 3056 12180 3108 12232
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4344 12223 4396 12232
rect 4068 12180 4120 12189
rect 4344 12189 4353 12223
rect 4353 12189 4387 12223
rect 4387 12189 4396 12223
rect 4344 12180 4396 12189
rect 5632 12223 5684 12232
rect 5632 12189 5641 12223
rect 5641 12189 5675 12223
rect 5675 12189 5684 12223
rect 5632 12180 5684 12189
rect 6552 12223 6604 12232
rect 6552 12189 6561 12223
rect 6561 12189 6595 12223
rect 6595 12189 6604 12223
rect 6552 12180 6604 12189
rect 7380 12223 7432 12232
rect 7380 12189 7389 12223
rect 7389 12189 7423 12223
rect 7423 12189 7432 12223
rect 7380 12180 7432 12189
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 8300 12180 8352 12232
rect 8484 12248 8536 12300
rect 9956 12384 10008 12436
rect 11888 12427 11940 12436
rect 11888 12393 11897 12427
rect 11897 12393 11931 12427
rect 11931 12393 11940 12427
rect 11888 12384 11940 12393
rect 14188 12384 14240 12436
rect 14832 12384 14884 12436
rect 9772 12316 9824 12368
rect 9956 12248 10008 12300
rect 12900 12248 12952 12300
rect 14648 12316 14700 12368
rect 9036 12180 9088 12232
rect 9312 12180 9364 12232
rect 9772 12223 9824 12232
rect 6184 12112 6236 12164
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 10692 12180 10744 12232
rect 11152 12180 11204 12232
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 7380 12044 7432 12096
rect 10140 12044 10192 12096
rect 11428 12112 11480 12164
rect 12440 12112 12492 12164
rect 11796 12044 11848 12096
rect 11980 12044 12032 12096
rect 12900 12044 12952 12096
rect 14464 12044 14516 12096
rect 5858 11942 5910 11994
rect 5922 11942 5974 11994
rect 5986 11942 6038 11994
rect 6050 11942 6102 11994
rect 10734 11942 10786 11994
rect 10798 11942 10850 11994
rect 10862 11942 10914 11994
rect 10926 11942 10978 11994
rect 1676 11883 1728 11892
rect 1676 11849 1685 11883
rect 1685 11849 1719 11883
rect 1719 11849 1728 11883
rect 1676 11840 1728 11849
rect 7012 11840 7064 11892
rect 8024 11883 8076 11892
rect 8024 11849 8033 11883
rect 8033 11849 8067 11883
rect 8067 11849 8076 11883
rect 8024 11840 8076 11849
rect 8484 11840 8536 11892
rect 6736 11815 6788 11824
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 3240 11704 3292 11756
rect 3792 11747 3844 11756
rect 3792 11713 3801 11747
rect 3801 11713 3835 11747
rect 3835 11713 3844 11747
rect 3792 11704 3844 11713
rect 4160 11704 4212 11756
rect 2964 11636 3016 11688
rect 5264 11704 5316 11756
rect 6736 11781 6745 11815
rect 6745 11781 6779 11815
rect 6779 11781 6788 11815
rect 6736 11772 6788 11781
rect 5632 11704 5684 11756
rect 6184 11704 6236 11756
rect 7012 11747 7064 11756
rect 7012 11713 7021 11747
rect 7021 11713 7055 11747
rect 7055 11713 7064 11747
rect 7012 11704 7064 11713
rect 7380 11704 7432 11756
rect 6460 11636 6512 11688
rect 6552 11636 6604 11688
rect 3056 11568 3108 11620
rect 3884 11500 3936 11552
rect 7748 11568 7800 11620
rect 7932 11704 7984 11756
rect 8116 11704 8168 11756
rect 9956 11840 10008 11892
rect 10140 11883 10192 11892
rect 10140 11849 10149 11883
rect 10149 11849 10183 11883
rect 10183 11849 10192 11883
rect 10140 11840 10192 11849
rect 11152 11840 11204 11892
rect 11336 11840 11388 11892
rect 9772 11772 9824 11824
rect 10692 11772 10744 11824
rect 12900 11815 12952 11824
rect 9036 11636 9088 11688
rect 11520 11704 11572 11756
rect 12900 11781 12909 11815
rect 12909 11781 12943 11815
rect 12943 11781 12952 11815
rect 12900 11772 12952 11781
rect 11888 11704 11940 11756
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 11152 11636 11204 11688
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 14832 11636 14884 11688
rect 11704 11568 11756 11620
rect 13820 11568 13872 11620
rect 7196 11500 7248 11552
rect 8024 11500 8076 11552
rect 9220 11500 9272 11552
rect 10324 11500 10376 11552
rect 10692 11500 10744 11552
rect 11980 11543 12032 11552
rect 11980 11509 11989 11543
rect 11989 11509 12023 11543
rect 12023 11509 12032 11543
rect 11980 11500 12032 11509
rect 12992 11500 13044 11552
rect 3420 11398 3472 11450
rect 3484 11398 3536 11450
rect 3548 11398 3600 11450
rect 3612 11398 3664 11450
rect 8296 11398 8348 11450
rect 8360 11398 8412 11450
rect 8424 11398 8476 11450
rect 8488 11398 8540 11450
rect 13172 11398 13224 11450
rect 13236 11398 13288 11450
rect 13300 11398 13352 11450
rect 13364 11398 13416 11450
rect 1952 11296 2004 11348
rect 3056 11296 3108 11348
rect 3148 11296 3200 11348
rect 5264 11339 5316 11348
rect 5264 11305 5273 11339
rect 5273 11305 5307 11339
rect 5307 11305 5316 11339
rect 5264 11296 5316 11305
rect 6460 11296 6512 11348
rect 7104 11296 7156 11348
rect 2044 11160 2096 11212
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 5632 11228 5684 11280
rect 7472 11228 7524 11280
rect 8116 11228 8168 11280
rect 9772 11228 9824 11280
rect 10600 11296 10652 11348
rect 11980 11296 12032 11348
rect 12716 11339 12768 11348
rect 12716 11305 12725 11339
rect 12725 11305 12759 11339
rect 12759 11305 12768 11339
rect 12716 11296 12768 11305
rect 12900 11296 12952 11348
rect 13912 11296 13964 11348
rect 14740 11296 14792 11348
rect 12808 11228 12860 11280
rect 3608 11092 3660 11144
rect 3792 11092 3844 11144
rect 4160 11092 4212 11144
rect 3148 11067 3200 11076
rect 3148 11033 3157 11067
rect 3157 11033 3191 11067
rect 3191 11033 3200 11067
rect 5724 11092 5776 11144
rect 7380 11160 7432 11212
rect 8668 11160 8720 11212
rect 11520 11160 11572 11212
rect 7840 11135 7892 11144
rect 3148 11024 3200 11033
rect 4988 11024 5040 11076
rect 5540 11067 5592 11076
rect 5540 11033 5549 11067
rect 5549 11033 5583 11067
rect 5583 11033 5592 11067
rect 5540 11024 5592 11033
rect 6276 11024 6328 11076
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 8852 11092 8904 11144
rect 11152 11135 11204 11144
rect 11152 11101 11161 11135
rect 11161 11101 11195 11135
rect 11195 11101 11204 11135
rect 12348 11160 12400 11212
rect 13084 11228 13136 11280
rect 13636 11228 13688 11280
rect 11888 11135 11940 11144
rect 11152 11092 11204 11101
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 12164 11092 12216 11144
rect 12900 11135 12952 11144
rect 12900 11101 12909 11135
rect 12909 11101 12943 11135
rect 12943 11101 12952 11135
rect 12900 11092 12952 11101
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 14556 11160 14608 11212
rect 12992 11092 13044 11101
rect 7472 11024 7524 11076
rect 7564 11024 7616 11076
rect 7932 11024 7984 11076
rect 4528 10956 4580 11008
rect 7104 10956 7156 11008
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 9312 11024 9364 11076
rect 10048 11067 10100 11076
rect 10048 11033 10057 11067
rect 10057 11033 10091 11067
rect 10091 11033 10100 11067
rect 10048 11024 10100 11033
rect 10232 11024 10284 11076
rect 10508 11024 10560 11076
rect 12440 11024 12492 11076
rect 13912 10956 13964 11008
rect 5858 10854 5910 10906
rect 5922 10854 5974 10906
rect 5986 10854 6038 10906
rect 6050 10854 6102 10906
rect 10734 10854 10786 10906
rect 10798 10854 10850 10906
rect 10862 10854 10914 10906
rect 10926 10854 10978 10906
rect 2044 10795 2096 10804
rect 2044 10761 2053 10795
rect 2053 10761 2087 10795
rect 2087 10761 2096 10795
rect 2044 10752 2096 10761
rect 3608 10795 3660 10804
rect 3608 10761 3617 10795
rect 3617 10761 3651 10795
rect 3651 10761 3660 10795
rect 3608 10752 3660 10761
rect 4896 10752 4948 10804
rect 4988 10752 5040 10804
rect 6552 10752 6604 10804
rect 6828 10752 6880 10804
rect 7288 10752 7340 10804
rect 9128 10752 9180 10804
rect 12072 10752 12124 10804
rect 2228 10659 2280 10668
rect 2228 10625 2237 10659
rect 2237 10625 2271 10659
rect 2271 10625 2280 10659
rect 2228 10616 2280 10625
rect 2504 10616 2556 10668
rect 2412 10548 2464 10600
rect 3240 10616 3292 10668
rect 5356 10684 5408 10736
rect 5540 10684 5592 10736
rect 4528 10659 4580 10668
rect 4528 10625 4537 10659
rect 4537 10625 4571 10659
rect 4571 10625 4580 10659
rect 4528 10616 4580 10625
rect 5724 10616 5776 10668
rect 9036 10684 9088 10736
rect 9772 10727 9824 10736
rect 7196 10659 7248 10668
rect 7196 10625 7205 10659
rect 7205 10625 7239 10659
rect 7239 10625 7248 10659
rect 7196 10616 7248 10625
rect 4620 10480 4672 10532
rect 6736 10480 6788 10532
rect 7840 10616 7892 10668
rect 7472 10591 7524 10600
rect 7472 10557 7481 10591
rect 7481 10557 7515 10591
rect 7515 10557 7524 10591
rect 7472 10548 7524 10557
rect 8944 10616 8996 10668
rect 9772 10693 9781 10727
rect 9781 10693 9815 10727
rect 9815 10693 9824 10727
rect 9772 10684 9824 10693
rect 10416 10684 10468 10736
rect 11980 10684 12032 10736
rect 9588 10616 9640 10668
rect 7564 10480 7616 10532
rect 7932 10480 7984 10532
rect 9864 10591 9916 10600
rect 9864 10557 9873 10591
rect 9873 10557 9907 10591
rect 9907 10557 9916 10591
rect 9864 10548 9916 10557
rect 10692 10659 10744 10668
rect 10692 10625 10701 10659
rect 10701 10625 10735 10659
rect 10735 10625 10744 10659
rect 10692 10616 10744 10625
rect 12072 10616 12124 10668
rect 12716 10616 12768 10668
rect 13084 10684 13136 10736
rect 13728 10659 13780 10668
rect 12624 10548 12676 10600
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 14648 10616 14700 10668
rect 13912 10548 13964 10600
rect 2688 10412 2740 10464
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 8116 10412 8168 10421
rect 8668 10412 8720 10464
rect 10600 10412 10652 10464
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 13084 10480 13136 10532
rect 14740 10480 14792 10532
rect 13728 10412 13780 10464
rect 3420 10310 3472 10362
rect 3484 10310 3536 10362
rect 3548 10310 3600 10362
rect 3612 10310 3664 10362
rect 8296 10310 8348 10362
rect 8360 10310 8412 10362
rect 8424 10310 8476 10362
rect 8488 10310 8540 10362
rect 13172 10310 13224 10362
rect 13236 10310 13288 10362
rect 13300 10310 13352 10362
rect 13364 10310 13416 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 3976 10208 4028 10260
rect 8852 10208 8904 10260
rect 10048 10208 10100 10260
rect 11888 10208 11940 10260
rect 12164 10208 12216 10260
rect 12992 10208 13044 10260
rect 2872 10140 2924 10192
rect 4436 10140 4488 10192
rect 12440 10183 12492 10192
rect 12440 10149 12449 10183
rect 12449 10149 12483 10183
rect 12483 10149 12492 10183
rect 12440 10140 12492 10149
rect 13084 10140 13136 10192
rect 14372 10140 14424 10192
rect 2688 10072 2740 10124
rect 4160 10047 4212 10056
rect 2228 9936 2280 9988
rect 2596 9979 2648 9988
rect 2596 9945 2605 9979
rect 2605 9945 2639 9979
rect 2639 9945 2648 9979
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 4896 10047 4948 10056
rect 4896 10013 4907 10047
rect 4907 10013 4948 10047
rect 4896 10004 4948 10013
rect 5632 10004 5684 10056
rect 7656 10004 7708 10056
rect 7748 10004 7800 10056
rect 7932 10047 7984 10056
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 8116 10047 8168 10056
rect 7932 10004 7984 10013
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 9312 10047 9364 10056
rect 9312 10013 9321 10047
rect 9321 10013 9355 10047
rect 9355 10013 9364 10047
rect 9312 10004 9364 10013
rect 2596 9936 2648 9945
rect 6552 9936 6604 9988
rect 4620 9868 4672 9920
rect 7012 9936 7064 9988
rect 7288 9936 7340 9988
rect 9036 9936 9088 9988
rect 9680 10072 9732 10124
rect 9864 10004 9916 10056
rect 11888 10072 11940 10124
rect 11060 10047 11112 10056
rect 11060 10013 11069 10047
rect 11069 10013 11103 10047
rect 11103 10013 11112 10047
rect 11060 10004 11112 10013
rect 11704 10004 11756 10056
rect 12164 10047 12216 10056
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 6920 9868 6972 9920
rect 7748 9868 7800 9920
rect 10232 9868 10284 9920
rect 11796 9936 11848 9988
rect 11888 9936 11940 9988
rect 12440 10004 12492 10056
rect 11244 9868 11296 9920
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 13728 10004 13780 10056
rect 13360 9936 13412 9988
rect 13084 9868 13136 9920
rect 5858 9766 5910 9818
rect 5922 9766 5974 9818
rect 5986 9766 6038 9818
rect 6050 9766 6102 9818
rect 10734 9766 10786 9818
rect 10798 9766 10850 9818
rect 10862 9766 10914 9818
rect 10926 9766 10978 9818
rect 2596 9664 2648 9716
rect 4160 9664 4212 9716
rect 6368 9664 6420 9716
rect 2688 9596 2740 9648
rect 2412 9460 2464 9512
rect 4988 9596 5040 9648
rect 9312 9664 9364 9716
rect 9588 9664 9640 9716
rect 10416 9664 10468 9716
rect 11152 9664 11204 9716
rect 11796 9664 11848 9716
rect 12440 9664 12492 9716
rect 12808 9664 12860 9716
rect 13268 9664 13320 9716
rect 2964 9392 3016 9444
rect 4436 9503 4488 9512
rect 4436 9469 4445 9503
rect 4445 9469 4479 9503
rect 4479 9469 4488 9503
rect 5632 9528 5684 9580
rect 5724 9528 5776 9580
rect 7012 9571 7064 9580
rect 7012 9537 7023 9571
rect 7023 9537 7064 9571
rect 5448 9503 5500 9512
rect 4436 9460 4488 9469
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 7012 9528 7064 9537
rect 7656 9528 7708 9580
rect 7932 9528 7984 9580
rect 7288 9460 7340 9512
rect 9128 9460 9180 9512
rect 9496 9460 9548 9512
rect 4712 9392 4764 9444
rect 9312 9392 9364 9444
rect 6368 9324 6420 9376
rect 7932 9324 7984 9376
rect 11888 9596 11940 9648
rect 9680 9460 9732 9512
rect 10324 9528 10376 9580
rect 11796 9571 11848 9580
rect 11796 9537 11805 9571
rect 11805 9537 11839 9571
rect 11839 9537 11848 9571
rect 11796 9528 11848 9537
rect 12808 9528 12860 9580
rect 13728 9528 13780 9580
rect 15108 9528 15160 9580
rect 10600 9460 10652 9512
rect 11704 9460 11756 9512
rect 12348 9460 12400 9512
rect 12900 9503 12952 9512
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 14280 9460 14332 9512
rect 14464 9460 14516 9512
rect 14832 9503 14884 9512
rect 14832 9469 14841 9503
rect 14841 9469 14875 9503
rect 14875 9469 14884 9503
rect 14832 9460 14884 9469
rect 13820 9392 13872 9444
rect 11060 9324 11112 9376
rect 12256 9324 12308 9376
rect 12992 9324 13044 9376
rect 3420 9222 3472 9274
rect 3484 9222 3536 9274
rect 3548 9222 3600 9274
rect 3612 9222 3664 9274
rect 8296 9222 8348 9274
rect 8360 9222 8412 9274
rect 8424 9222 8476 9274
rect 8488 9222 8540 9274
rect 13172 9222 13224 9274
rect 13236 9222 13288 9274
rect 13300 9222 13352 9274
rect 13364 9222 13416 9274
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 5448 9120 5500 9172
rect 6368 9163 6420 9172
rect 6368 9129 6377 9163
rect 6377 9129 6411 9163
rect 6411 9129 6420 9163
rect 6368 9120 6420 9129
rect 7012 9120 7064 9172
rect 8116 9120 8168 9172
rect 8760 9120 8812 9172
rect 9036 9120 9088 9172
rect 9312 9163 9364 9172
rect 9312 9129 9321 9163
rect 9321 9129 9355 9163
rect 9355 9129 9364 9163
rect 9312 9120 9364 9129
rect 11428 9120 11480 9172
rect 12808 9163 12860 9172
rect 11060 9052 11112 9104
rect 3976 8984 4028 9036
rect 7380 8984 7432 9036
rect 7472 8984 7524 9036
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 3792 8959 3844 8968
rect 1860 8848 1912 8900
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 4436 8916 4488 8968
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4988 8959 5040 8968
rect 4712 8916 4764 8925
rect 4988 8925 4997 8959
rect 4997 8925 5031 8959
rect 5031 8925 5040 8959
rect 4988 8916 5040 8925
rect 6920 8916 6972 8968
rect 3976 8823 4028 8832
rect 3976 8789 3985 8823
rect 3985 8789 4019 8823
rect 4019 8789 4028 8823
rect 3976 8780 4028 8789
rect 4068 8780 4120 8832
rect 6552 8848 6604 8900
rect 7288 8916 7340 8968
rect 12808 9129 12817 9163
rect 12817 9129 12851 9163
rect 12851 9129 12860 9163
rect 12808 9120 12860 9129
rect 14464 9163 14516 9172
rect 14464 9129 14473 9163
rect 14473 9129 14507 9163
rect 14507 9129 14516 9163
rect 14464 9120 14516 9129
rect 12440 9052 12492 9104
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 8944 8891 8996 8900
rect 8944 8857 8953 8891
rect 8953 8857 8987 8891
rect 8987 8857 8996 8891
rect 8944 8848 8996 8857
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 7472 8780 7524 8832
rect 9864 8916 9916 8968
rect 11428 8916 11480 8968
rect 11612 8959 11664 8968
rect 11612 8925 11621 8959
rect 11621 8925 11655 8959
rect 11655 8925 11664 8959
rect 11612 8916 11664 8925
rect 13820 8916 13872 8968
rect 14372 8916 14424 8968
rect 10416 8848 10468 8900
rect 9588 8780 9640 8832
rect 15016 8848 15068 8900
rect 11980 8823 12032 8832
rect 11980 8789 11989 8823
rect 11989 8789 12023 8823
rect 12023 8789 12032 8823
rect 11980 8780 12032 8789
rect 5858 8678 5910 8730
rect 5922 8678 5974 8730
rect 5986 8678 6038 8730
rect 6050 8678 6102 8730
rect 10734 8678 10786 8730
rect 10798 8678 10850 8730
rect 10862 8678 10914 8730
rect 10926 8678 10978 8730
rect 5448 8576 5500 8628
rect 3148 8508 3200 8560
rect 2780 8440 2832 8492
rect 4068 8508 4120 8560
rect 2320 8415 2372 8424
rect 2320 8381 2329 8415
rect 2329 8381 2363 8415
rect 2363 8381 2372 8415
rect 2320 8372 2372 8381
rect 2872 8347 2924 8356
rect 2872 8313 2881 8347
rect 2881 8313 2915 8347
rect 2915 8313 2924 8347
rect 2872 8304 2924 8313
rect 3884 8483 3936 8492
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 6920 8508 6972 8560
rect 3884 8440 3936 8449
rect 6368 8440 6420 8492
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 9220 8508 9272 8560
rect 8668 8440 8720 8492
rect 8944 8440 8996 8492
rect 10508 8576 10560 8628
rect 11244 8576 11296 8628
rect 13728 8576 13780 8628
rect 14464 8576 14516 8628
rect 15200 8576 15252 8628
rect 11060 8508 11112 8560
rect 12992 8508 13044 8560
rect 9588 8483 9640 8492
rect 8760 8372 8812 8424
rect 9588 8449 9597 8483
rect 9597 8449 9631 8483
rect 9631 8449 9640 8483
rect 10416 8483 10468 8492
rect 9588 8440 9640 8449
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 11520 8440 11572 8492
rect 9496 8415 9548 8424
rect 5908 8304 5960 8356
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 11060 8372 11112 8424
rect 11612 8372 11664 8424
rect 11888 8372 11940 8424
rect 12900 8440 12952 8492
rect 13544 8440 13596 8492
rect 12808 8372 12860 8424
rect 13452 8372 13504 8424
rect 14280 8440 14332 8492
rect 14004 8415 14056 8424
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 1860 8236 1912 8288
rect 3148 8236 3200 8288
rect 5172 8279 5224 8288
rect 5172 8245 5181 8279
rect 5181 8245 5215 8279
rect 5215 8245 5224 8279
rect 5172 8236 5224 8245
rect 9312 8304 9364 8356
rect 7380 8279 7432 8288
rect 7380 8245 7389 8279
rect 7389 8245 7423 8279
rect 7423 8245 7432 8279
rect 7380 8236 7432 8245
rect 9864 8304 9916 8356
rect 14556 8304 14608 8356
rect 14832 8304 14884 8356
rect 9956 8236 10008 8288
rect 10692 8236 10744 8288
rect 12716 8236 12768 8288
rect 12900 8279 12952 8288
rect 12900 8245 12909 8279
rect 12909 8245 12943 8279
rect 12943 8245 12952 8279
rect 12900 8236 12952 8245
rect 3420 8134 3472 8186
rect 3484 8134 3536 8186
rect 3548 8134 3600 8186
rect 3612 8134 3664 8186
rect 8296 8134 8348 8186
rect 8360 8134 8412 8186
rect 8424 8134 8476 8186
rect 8488 8134 8540 8186
rect 13172 8134 13224 8186
rect 13236 8134 13288 8186
rect 13300 8134 13352 8186
rect 13364 8134 13416 8186
rect 2320 8032 2372 8084
rect 10508 8032 10560 8084
rect 10600 8032 10652 8084
rect 3148 7939 3200 7948
rect 3148 7905 3157 7939
rect 3157 7905 3191 7939
rect 3191 7905 3200 7939
rect 3148 7896 3200 7905
rect 3700 7964 3752 8016
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 2688 7828 2740 7880
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 5172 7896 5224 7948
rect 5724 7964 5776 8016
rect 10416 7964 10468 8016
rect 13820 7964 13872 8016
rect 6920 7896 6972 7948
rect 6736 7871 6788 7880
rect 2136 7692 2188 7744
rect 5540 7760 5592 7812
rect 5908 7760 5960 7812
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 6276 7760 6328 7812
rect 6460 7803 6512 7812
rect 6460 7769 6469 7803
rect 6469 7769 6503 7803
rect 6503 7769 6512 7803
rect 6460 7760 6512 7769
rect 6828 7760 6880 7812
rect 7564 7828 7616 7880
rect 11704 7896 11756 7948
rect 9588 7871 9640 7880
rect 9588 7837 9597 7871
rect 9597 7837 9631 7871
rect 9631 7837 9640 7871
rect 9588 7828 9640 7837
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 11060 7871 11112 7880
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 11888 7828 11940 7880
rect 9496 7803 9548 7812
rect 9496 7769 9505 7803
rect 9505 7769 9539 7803
rect 9539 7769 9548 7803
rect 9496 7760 9548 7769
rect 10048 7760 10100 7812
rect 11612 7760 11664 7812
rect 12716 7828 12768 7880
rect 12532 7760 12584 7812
rect 13544 7828 13596 7880
rect 14280 7828 14332 7880
rect 13728 7760 13780 7812
rect 7472 7692 7524 7744
rect 11336 7692 11388 7744
rect 11704 7692 11756 7744
rect 12992 7735 13044 7744
rect 12992 7701 13001 7735
rect 13001 7701 13035 7735
rect 13035 7701 13044 7735
rect 12992 7692 13044 7701
rect 5858 7590 5910 7642
rect 5922 7590 5974 7642
rect 5986 7590 6038 7642
rect 6050 7590 6102 7642
rect 10734 7590 10786 7642
rect 10798 7590 10850 7642
rect 10862 7590 10914 7642
rect 10926 7590 10978 7642
rect 6920 7531 6972 7540
rect 3148 7420 3200 7472
rect 2872 7395 2924 7404
rect 2872 7361 2881 7395
rect 2881 7361 2915 7395
rect 2915 7361 2924 7395
rect 2872 7352 2924 7361
rect 3700 7395 3752 7404
rect 3700 7361 3709 7395
rect 3709 7361 3743 7395
rect 3743 7361 3752 7395
rect 3700 7352 3752 7361
rect 5172 7420 5224 7472
rect 6920 7497 6929 7531
rect 6929 7497 6963 7531
rect 6963 7497 6972 7531
rect 6920 7488 6972 7497
rect 10048 7488 10100 7540
rect 10416 7488 10468 7540
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 3884 7284 3936 7336
rect 7012 7352 7064 7404
rect 7840 7420 7892 7472
rect 5540 7284 5592 7336
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7564 7395 7616 7404
rect 7564 7361 7573 7395
rect 7573 7361 7607 7395
rect 7607 7361 7616 7395
rect 7564 7352 7616 7361
rect 11888 7420 11940 7472
rect 12532 7463 12584 7472
rect 12532 7429 12541 7463
rect 12541 7429 12575 7463
rect 12575 7429 12584 7463
rect 12532 7420 12584 7429
rect 12900 7420 12952 7472
rect 13544 7488 13596 7540
rect 9864 7352 9916 7404
rect 10232 7352 10284 7404
rect 11152 7352 11204 7404
rect 11796 7352 11848 7404
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 7288 7284 7340 7293
rect 10968 7284 11020 7336
rect 11980 7284 12032 7336
rect 13084 7352 13136 7404
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 13820 7284 13872 7336
rect 13912 7284 13964 7336
rect 14372 7327 14424 7336
rect 14372 7293 14381 7327
rect 14381 7293 14415 7327
rect 14415 7293 14424 7327
rect 14372 7284 14424 7293
rect 3240 7148 3292 7200
rect 5264 7148 5316 7200
rect 5724 7148 5776 7200
rect 12532 7216 12584 7268
rect 7472 7148 7524 7200
rect 8944 7148 8996 7200
rect 10140 7148 10192 7200
rect 11060 7148 11112 7200
rect 11152 7148 11204 7200
rect 12072 7148 12124 7200
rect 12256 7191 12308 7200
rect 12256 7157 12265 7191
rect 12265 7157 12299 7191
rect 12299 7157 12308 7191
rect 12256 7148 12308 7157
rect 12440 7148 12492 7200
rect 12808 7148 12860 7200
rect 13820 7148 13872 7200
rect 3420 7046 3472 7098
rect 3484 7046 3536 7098
rect 3548 7046 3600 7098
rect 3612 7046 3664 7098
rect 8296 7046 8348 7098
rect 8360 7046 8412 7098
rect 8424 7046 8476 7098
rect 8488 7046 8540 7098
rect 13172 7046 13224 7098
rect 13236 7046 13288 7098
rect 13300 7046 13352 7098
rect 13364 7046 13416 7098
rect 2872 6944 2924 6996
rect 8852 6944 8904 6996
rect 10600 6944 10652 6996
rect 10968 6987 11020 6996
rect 10968 6953 10977 6987
rect 10977 6953 11011 6987
rect 11011 6953 11020 6987
rect 10968 6944 11020 6953
rect 11060 6944 11112 6996
rect 11612 6944 11664 6996
rect 11980 6944 12032 6996
rect 12348 6944 12400 6996
rect 12808 6944 12860 6996
rect 1584 6740 1636 6792
rect 2136 6808 2188 6860
rect 4436 6808 4488 6860
rect 5264 6808 5316 6860
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4068 6783 4120 6792
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 5172 6783 5224 6792
rect 3240 6672 3292 6724
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 5172 6740 5224 6749
rect 6276 6740 6328 6792
rect 7288 6808 7340 6860
rect 7656 6851 7708 6860
rect 7656 6817 7665 6851
rect 7665 6817 7699 6851
rect 7699 6817 7708 6851
rect 7656 6808 7708 6817
rect 6828 6783 6880 6792
rect 1584 6604 1636 6656
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 3056 6604 3108 6656
rect 4988 6604 5040 6656
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 10416 6808 10468 6860
rect 7840 6740 7892 6792
rect 7932 6740 7984 6792
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 8668 6740 8720 6792
rect 6736 6672 6788 6724
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 7564 6604 7616 6656
rect 8484 6604 8536 6656
rect 9864 6740 9916 6792
rect 10232 6672 10284 6724
rect 12256 6783 12308 6792
rect 12256 6749 12265 6783
rect 12265 6749 12299 6783
rect 12299 6749 12308 6783
rect 12256 6740 12308 6749
rect 12900 6740 12952 6792
rect 13728 6808 13780 6860
rect 14372 6851 14424 6860
rect 14372 6817 14381 6851
rect 14381 6817 14415 6851
rect 14415 6817 14424 6851
rect 14372 6808 14424 6817
rect 13636 6740 13688 6792
rect 12992 6672 13044 6724
rect 12164 6604 12216 6656
rect 14648 6604 14700 6656
rect 5858 6502 5910 6554
rect 5922 6502 5974 6554
rect 5986 6502 6038 6554
rect 6050 6502 6102 6554
rect 10734 6502 10786 6554
rect 10798 6502 10850 6554
rect 10862 6502 10914 6554
rect 10926 6502 10978 6554
rect 1676 6400 1728 6452
rect 4068 6400 4120 6452
rect 4436 6443 4488 6452
rect 4436 6409 4445 6443
rect 4445 6409 4479 6443
rect 4479 6409 4488 6443
rect 4436 6400 4488 6409
rect 3240 6332 3292 6384
rect 1584 6196 1636 6248
rect 4896 6332 4948 6384
rect 6368 6332 6420 6384
rect 6828 6332 6880 6384
rect 7104 6375 7156 6384
rect 7104 6341 7113 6375
rect 7113 6341 7147 6375
rect 7147 6341 7156 6375
rect 8852 6400 8904 6452
rect 9588 6443 9640 6452
rect 9588 6409 9597 6443
rect 9597 6409 9631 6443
rect 9631 6409 9640 6443
rect 9588 6400 9640 6409
rect 11704 6400 11756 6452
rect 11796 6400 11848 6452
rect 14280 6400 14332 6452
rect 7104 6332 7156 6341
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 6276 6264 6328 6316
rect 7196 6264 7248 6316
rect 4988 6239 5040 6248
rect 4988 6205 4997 6239
rect 4997 6205 5031 6239
rect 5031 6205 5040 6239
rect 4988 6196 5040 6205
rect 8116 6332 8168 6384
rect 8484 6375 8536 6384
rect 8484 6341 8493 6375
rect 8493 6341 8527 6375
rect 8527 6341 8536 6375
rect 8484 6332 8536 6341
rect 8576 6332 8628 6384
rect 9312 6332 9364 6384
rect 11060 6332 11112 6384
rect 11336 6332 11388 6384
rect 9956 6264 10008 6316
rect 10784 6307 10836 6316
rect 10784 6273 10793 6307
rect 10793 6273 10827 6307
rect 10827 6273 10836 6307
rect 10784 6264 10836 6273
rect 11796 6307 11848 6316
rect 11796 6273 11805 6307
rect 11805 6273 11839 6307
rect 11839 6273 11848 6307
rect 11796 6264 11848 6273
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 11980 6264 12032 6273
rect 12808 6307 12860 6316
rect 12808 6273 12817 6307
rect 12817 6273 12851 6307
rect 12851 6273 12860 6307
rect 12808 6264 12860 6273
rect 8024 6196 8076 6248
rect 9588 6196 9640 6248
rect 11152 6196 11204 6248
rect 11612 6196 11664 6248
rect 2596 6128 2648 6180
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 3240 6128 3292 6180
rect 6368 6128 6420 6180
rect 9128 6128 9180 6180
rect 9312 6171 9364 6180
rect 9312 6137 9321 6171
rect 9321 6137 9355 6171
rect 9355 6137 9364 6171
rect 9312 6128 9364 6137
rect 9496 6128 9548 6180
rect 10140 6128 10192 6180
rect 10324 6128 10376 6180
rect 12992 6307 13044 6316
rect 12992 6273 13001 6307
rect 13001 6273 13035 6307
rect 13035 6273 13044 6307
rect 12992 6264 13044 6273
rect 13820 6307 13872 6316
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 13820 6264 13872 6273
rect 14556 6196 14608 6248
rect 6000 6060 6052 6112
rect 7104 6060 7156 6112
rect 8944 6060 8996 6112
rect 10876 6060 10928 6112
rect 10968 6103 11020 6112
rect 10968 6069 10977 6103
rect 10977 6069 11011 6103
rect 11011 6069 11020 6103
rect 12992 6128 13044 6180
rect 12164 6103 12216 6112
rect 10968 6060 11020 6069
rect 12164 6069 12173 6103
rect 12173 6069 12207 6103
rect 12207 6069 12216 6103
rect 12164 6060 12216 6069
rect 12256 6060 12308 6112
rect 14832 6060 14884 6112
rect 3420 5958 3472 6010
rect 3484 5958 3536 6010
rect 3548 5958 3600 6010
rect 3612 5958 3664 6010
rect 8296 5958 8348 6010
rect 8360 5958 8412 6010
rect 8424 5958 8476 6010
rect 8488 5958 8540 6010
rect 13172 5958 13224 6010
rect 13236 5958 13288 6010
rect 13300 5958 13352 6010
rect 13364 5958 13416 6010
rect 2044 5856 2096 5908
rect 3240 5831 3292 5840
rect 3240 5797 3249 5831
rect 3249 5797 3283 5831
rect 3283 5797 3292 5831
rect 3240 5788 3292 5797
rect 3976 5763 4028 5772
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 7380 5788 7432 5840
rect 9220 5856 9272 5908
rect 3976 5720 4028 5729
rect 2136 5652 2188 5704
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 2320 5584 2372 5636
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 5356 5652 5408 5704
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 8024 5695 8076 5704
rect 6920 5652 6972 5661
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8392 5695 8444 5704
rect 8116 5652 8168 5661
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 9864 5788 9916 5840
rect 10048 5831 10100 5840
rect 10048 5797 10057 5831
rect 10057 5797 10091 5831
rect 10091 5797 10100 5831
rect 10048 5788 10100 5797
rect 12808 5856 12860 5908
rect 14464 5856 14516 5908
rect 11980 5788 12032 5840
rect 1584 5516 1636 5568
rect 2596 5559 2648 5568
rect 2596 5525 2605 5559
rect 2605 5525 2639 5559
rect 2639 5525 2648 5559
rect 2596 5516 2648 5525
rect 6736 5584 6788 5636
rect 7104 5627 7156 5636
rect 7104 5593 7113 5627
rect 7113 5593 7147 5627
rect 7147 5593 7156 5627
rect 7104 5584 7156 5593
rect 10600 5652 10652 5704
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 10968 5695 11020 5704
rect 10968 5661 10977 5695
rect 10977 5661 11011 5695
rect 11011 5661 11020 5695
rect 10968 5652 11020 5661
rect 14004 5788 14056 5840
rect 14280 5788 14332 5840
rect 14372 5763 14424 5772
rect 14372 5729 14381 5763
rect 14381 5729 14415 5763
rect 14415 5729 14424 5763
rect 14372 5720 14424 5729
rect 14556 5720 14608 5772
rect 9772 5584 9824 5636
rect 10508 5584 10560 5636
rect 12348 5652 12400 5704
rect 12808 5652 12860 5704
rect 13452 5652 13504 5704
rect 13820 5652 13872 5704
rect 14556 5584 14608 5636
rect 14832 5584 14884 5636
rect 14924 5584 14976 5636
rect 5632 5516 5684 5568
rect 7840 5559 7892 5568
rect 7840 5525 7849 5559
rect 7849 5525 7883 5559
rect 7883 5525 7892 5559
rect 7840 5516 7892 5525
rect 8208 5516 8260 5568
rect 9680 5516 9732 5568
rect 10140 5516 10192 5568
rect 10324 5516 10376 5568
rect 11796 5516 11848 5568
rect 12808 5559 12860 5568
rect 12808 5525 12817 5559
rect 12817 5525 12851 5559
rect 12851 5525 12860 5559
rect 12808 5516 12860 5525
rect 14004 5516 14056 5568
rect 5858 5414 5910 5466
rect 5922 5414 5974 5466
rect 5986 5414 6038 5466
rect 6050 5414 6102 5466
rect 10734 5414 10786 5466
rect 10798 5414 10850 5466
rect 10862 5414 10914 5466
rect 10926 5414 10978 5466
rect 2872 5312 2924 5364
rect 3148 5312 3200 5364
rect 4620 5244 4672 5296
rect 6920 5312 6972 5364
rect 9772 5312 9824 5364
rect 9864 5312 9916 5364
rect 10508 5355 10560 5364
rect 10508 5321 10517 5355
rect 10517 5321 10551 5355
rect 10551 5321 10560 5355
rect 10508 5312 10560 5321
rect 11612 5355 11664 5364
rect 11612 5321 11621 5355
rect 11621 5321 11655 5355
rect 11655 5321 11664 5355
rect 11612 5312 11664 5321
rect 12992 5312 13044 5364
rect 14188 5355 14240 5364
rect 14188 5321 14197 5355
rect 14197 5321 14231 5355
rect 14231 5321 14240 5355
rect 14188 5312 14240 5321
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 3148 5176 3200 5228
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 4344 5176 4396 5228
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 4988 5219 5040 5228
rect 4988 5185 4997 5219
rect 4997 5185 5031 5219
rect 5031 5185 5040 5219
rect 5264 5219 5316 5228
rect 4988 5176 5040 5185
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 7012 5176 7064 5228
rect 5172 5151 5224 5160
rect 5172 5117 5181 5151
rect 5181 5117 5215 5151
rect 5215 5117 5224 5151
rect 5172 5108 5224 5117
rect 6552 5108 6604 5160
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 8760 5219 8812 5228
rect 8760 5185 8769 5219
rect 8769 5185 8803 5219
rect 8803 5185 8812 5219
rect 8760 5176 8812 5185
rect 8944 5176 8996 5228
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 9404 5176 9456 5228
rect 11520 5244 11572 5296
rect 13912 5244 13964 5296
rect 10048 5219 10100 5228
rect 10048 5185 10057 5219
rect 10057 5185 10091 5219
rect 10091 5185 10100 5219
rect 10048 5176 10100 5185
rect 10140 5219 10192 5228
rect 10140 5185 10149 5219
rect 10149 5185 10183 5219
rect 10183 5185 10192 5219
rect 10140 5176 10192 5185
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 11796 5219 11848 5228
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 11980 5219 12032 5228
rect 11796 5176 11848 5185
rect 11980 5185 11989 5219
rect 11989 5185 12023 5219
rect 12023 5185 12032 5219
rect 11980 5176 12032 5185
rect 12164 5176 12216 5228
rect 12440 5176 12492 5228
rect 12992 5219 13044 5228
rect 12992 5185 13001 5219
rect 13001 5185 13035 5219
rect 13035 5185 13044 5219
rect 12992 5176 13044 5185
rect 13452 5176 13504 5228
rect 14280 5219 14332 5228
rect 14280 5185 14289 5219
rect 14289 5185 14323 5219
rect 14323 5185 14332 5219
rect 14280 5176 14332 5185
rect 15016 5219 15068 5228
rect 15016 5185 15025 5219
rect 15025 5185 15059 5219
rect 15059 5185 15068 5219
rect 15016 5176 15068 5185
rect 10600 5108 10652 5160
rect 11520 5108 11572 5160
rect 13636 5108 13688 5160
rect 4068 5040 4120 5092
rect 4252 5040 4304 5092
rect 7564 5040 7616 5092
rect 8116 5040 8168 5092
rect 8944 5040 8996 5092
rect 9404 5040 9456 5092
rect 10416 5040 10468 5092
rect 14464 5040 14516 5092
rect 3792 4972 3844 5024
rect 4712 4972 4764 5024
rect 9128 4972 9180 5024
rect 9312 5015 9364 5024
rect 9312 4981 9321 5015
rect 9321 4981 9355 5015
rect 9355 4981 9364 5015
rect 9312 4972 9364 4981
rect 12440 4972 12492 5024
rect 14188 4972 14240 5024
rect 3420 4870 3472 4922
rect 3484 4870 3536 4922
rect 3548 4870 3600 4922
rect 3612 4870 3664 4922
rect 8296 4870 8348 4922
rect 8360 4870 8412 4922
rect 8424 4870 8476 4922
rect 8488 4870 8540 4922
rect 13172 4870 13224 4922
rect 13236 4870 13288 4922
rect 13300 4870 13352 4922
rect 13364 4870 13416 4922
rect 2044 4700 2096 4752
rect 3976 4768 4028 4820
rect 8024 4768 8076 4820
rect 10324 4768 10376 4820
rect 11060 4768 11112 4820
rect 12992 4768 13044 4820
rect 4068 4700 4120 4752
rect 6276 4700 6328 4752
rect 8852 4700 8904 4752
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 2412 4564 2464 4616
rect 4160 4632 4212 4684
rect 4344 4675 4396 4684
rect 4344 4641 4353 4675
rect 4353 4641 4387 4675
rect 4387 4641 4396 4675
rect 4344 4632 4396 4641
rect 3056 4607 3108 4616
rect 2136 4496 2188 4548
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 7012 4632 7064 4684
rect 7840 4632 7892 4684
rect 8668 4632 8720 4684
rect 9680 4632 9732 4684
rect 10508 4632 10560 4684
rect 5724 4564 5776 4616
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7380 4607 7432 4616
rect 7380 4573 7389 4607
rect 7389 4573 7423 4607
rect 7423 4573 7432 4607
rect 7380 4564 7432 4573
rect 8116 4564 8168 4616
rect 9220 4564 9272 4616
rect 9588 4607 9640 4616
rect 9588 4573 9600 4607
rect 9600 4573 9634 4607
rect 9634 4573 9640 4607
rect 9588 4564 9640 4573
rect 11060 4564 11112 4616
rect 8944 4496 8996 4548
rect 9680 4496 9732 4548
rect 10232 4496 10284 4548
rect 11888 4700 11940 4752
rect 12532 4700 12584 4752
rect 11796 4632 11848 4684
rect 11520 4607 11572 4616
rect 11520 4573 11529 4607
rect 11529 4573 11563 4607
rect 11563 4573 11572 4607
rect 11520 4564 11572 4573
rect 11888 4607 11940 4616
rect 11888 4573 11897 4607
rect 11897 4573 11931 4607
rect 11931 4573 11940 4607
rect 12716 4632 12768 4684
rect 14188 4700 14240 4752
rect 14464 4675 14516 4684
rect 13084 4607 13136 4616
rect 11888 4564 11940 4573
rect 13084 4573 13093 4607
rect 13093 4573 13127 4607
rect 13127 4573 13136 4607
rect 13084 4564 13136 4573
rect 13268 4607 13320 4616
rect 13268 4573 13277 4607
rect 13277 4573 13311 4607
rect 13311 4573 13320 4607
rect 13268 4564 13320 4573
rect 13360 4607 13412 4616
rect 13360 4573 13395 4607
rect 13395 4573 13412 4607
rect 13544 4607 13596 4636
rect 13544 4584 13553 4607
rect 13553 4584 13587 4607
rect 13587 4584 13596 4607
rect 14464 4641 14473 4675
rect 14473 4641 14507 4675
rect 14507 4641 14516 4675
rect 14464 4632 14516 4641
rect 14648 4700 14700 4752
rect 13360 4564 13412 4573
rect 13728 4564 13780 4616
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 11612 4539 11664 4548
rect 2964 4471 3016 4480
rect 2964 4437 2973 4471
rect 2973 4437 3007 4471
rect 3007 4437 3016 4471
rect 2964 4428 3016 4437
rect 4344 4428 4396 4480
rect 7104 4471 7156 4480
rect 7104 4437 7113 4471
rect 7113 4437 7147 4471
rect 7147 4437 7156 4471
rect 7104 4428 7156 4437
rect 8208 4428 8260 4480
rect 9404 4428 9456 4480
rect 10140 4428 10192 4480
rect 11060 4428 11112 4480
rect 11612 4505 11621 4539
rect 11621 4505 11655 4539
rect 11655 4505 11664 4539
rect 11612 4496 11664 4505
rect 12808 4496 12860 4548
rect 12532 4428 12584 4480
rect 13912 4496 13964 4548
rect 13084 4428 13136 4480
rect 5858 4326 5910 4378
rect 5922 4326 5974 4378
rect 5986 4326 6038 4378
rect 6050 4326 6102 4378
rect 10734 4326 10786 4378
rect 10798 4326 10850 4378
rect 10862 4326 10914 4378
rect 10926 4326 10978 4378
rect 2964 4224 3016 4276
rect 4712 4224 4764 4276
rect 6368 4224 6420 4276
rect 8944 4267 8996 4276
rect 8944 4233 8953 4267
rect 8953 4233 8987 4267
rect 8987 4233 8996 4267
rect 8944 4224 8996 4233
rect 9588 4224 9640 4276
rect 12716 4224 12768 4276
rect 12900 4224 12952 4276
rect 14464 4267 14516 4276
rect 14464 4233 14473 4267
rect 14473 4233 14507 4267
rect 14507 4233 14516 4267
rect 14464 4224 14516 4233
rect 4344 4199 4396 4208
rect 4344 4165 4353 4199
rect 4353 4165 4387 4199
rect 4387 4165 4396 4199
rect 4344 4156 4396 4165
rect 6184 4156 6236 4208
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 3976 4131 4028 4140
rect 2964 4020 3016 4072
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 7012 4131 7064 4140
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 7012 4088 7064 4097
rect 7104 4088 7156 4140
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 8668 4088 8720 4140
rect 9312 4156 9364 4208
rect 12808 4156 12860 4208
rect 12992 4156 13044 4208
rect 9128 4088 9180 4140
rect 9220 4088 9272 4140
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 11704 4131 11756 4140
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 11980 4088 12032 4140
rect 5724 3952 5776 4004
rect 2964 3884 3016 3936
rect 5080 3884 5132 3936
rect 7288 3952 7340 4004
rect 9404 3952 9456 4004
rect 11888 4020 11940 4072
rect 12624 4088 12676 4140
rect 13360 4088 13412 4140
rect 14188 4131 14240 4140
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 14188 4088 14240 4097
rect 14280 4131 14332 4140
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 14648 4088 14700 4140
rect 13544 4020 13596 4072
rect 11980 3952 12032 4004
rect 13452 3952 13504 4004
rect 13912 3952 13964 4004
rect 7472 3884 7524 3936
rect 9588 3927 9640 3936
rect 9588 3893 9597 3927
rect 9597 3893 9631 3927
rect 9631 3893 9640 3927
rect 9588 3884 9640 3893
rect 11244 3884 11296 3936
rect 3420 3782 3472 3834
rect 3484 3782 3536 3834
rect 3548 3782 3600 3834
rect 3612 3782 3664 3834
rect 8296 3782 8348 3834
rect 8360 3782 8412 3834
rect 8424 3782 8476 3834
rect 8488 3782 8540 3834
rect 13172 3782 13224 3834
rect 13236 3782 13288 3834
rect 13300 3782 13352 3834
rect 13364 3782 13416 3834
rect 12624 3680 12676 3732
rect 14096 3723 14148 3732
rect 14096 3689 14105 3723
rect 14105 3689 14139 3723
rect 14139 3689 14148 3723
rect 14096 3680 14148 3689
rect 5080 3655 5132 3664
rect 5080 3621 5089 3655
rect 5089 3621 5123 3655
rect 5123 3621 5132 3655
rect 5080 3612 5132 3621
rect 6460 3612 6512 3664
rect 2780 3544 2832 3596
rect 4988 3544 5040 3596
rect 6920 3544 6972 3596
rect 7656 3544 7708 3596
rect 8668 3612 8720 3664
rect 12716 3612 12768 3664
rect 9588 3587 9640 3596
rect 3240 3519 3292 3528
rect 3240 3485 3249 3519
rect 3249 3485 3283 3519
rect 3283 3485 3292 3519
rect 3240 3476 3292 3485
rect 3700 3476 3752 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 3608 3408 3660 3460
rect 4160 3408 4212 3460
rect 5356 3476 5408 3528
rect 6368 3476 6420 3528
rect 6460 3476 6512 3528
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7196 3519 7248 3528
rect 7012 3476 7064 3485
rect 7196 3485 7205 3519
rect 7205 3485 7239 3519
rect 7239 3485 7248 3519
rect 7196 3476 7248 3485
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7472 3519 7524 3528
rect 7288 3476 7340 3485
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 2964 3340 3016 3392
rect 3792 3340 3844 3392
rect 7656 3408 7708 3460
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 8760 3476 8812 3528
rect 7104 3340 7156 3392
rect 7840 3340 7892 3392
rect 8024 3383 8076 3392
rect 8024 3349 8033 3383
rect 8033 3349 8067 3383
rect 8067 3349 8076 3383
rect 8024 3340 8076 3349
rect 9588 3553 9597 3587
rect 9597 3553 9631 3587
rect 9631 3553 9640 3587
rect 9588 3544 9640 3553
rect 9864 3544 9916 3596
rect 9680 3476 9732 3528
rect 12900 3544 12952 3596
rect 14464 3587 14516 3596
rect 14464 3553 14473 3587
rect 14473 3553 14507 3587
rect 14507 3553 14516 3587
rect 14464 3544 14516 3553
rect 10140 3476 10192 3528
rect 11060 3519 11112 3528
rect 11060 3485 11069 3519
rect 11069 3485 11103 3519
rect 11103 3485 11112 3519
rect 11060 3476 11112 3485
rect 11244 3519 11296 3528
rect 11244 3485 11253 3519
rect 11253 3485 11287 3519
rect 11287 3485 11296 3519
rect 11244 3476 11296 3485
rect 11888 3519 11940 3528
rect 11888 3485 11897 3519
rect 11897 3485 11931 3519
rect 11931 3485 11940 3519
rect 11888 3476 11940 3485
rect 9864 3408 9916 3460
rect 11152 3451 11204 3460
rect 11152 3417 11161 3451
rect 11161 3417 11195 3451
rect 11195 3417 11204 3451
rect 11152 3408 11204 3417
rect 12256 3519 12308 3528
rect 12256 3485 12265 3519
rect 12265 3485 12299 3519
rect 12299 3485 12308 3519
rect 12256 3476 12308 3485
rect 14004 3476 14056 3528
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 14648 3476 14700 3528
rect 13544 3451 13596 3460
rect 13544 3417 13553 3451
rect 13553 3417 13587 3451
rect 13587 3417 13596 3451
rect 13544 3408 13596 3417
rect 11796 3340 11848 3392
rect 13636 3340 13688 3392
rect 5858 3238 5910 3290
rect 5922 3238 5974 3290
rect 5986 3238 6038 3290
rect 6050 3238 6102 3290
rect 10734 3238 10786 3290
rect 10798 3238 10850 3290
rect 10862 3238 10914 3290
rect 10926 3238 10978 3290
rect 1400 2975 1452 2984
rect 1400 2941 1409 2975
rect 1409 2941 1443 2975
rect 1443 2941 1452 2975
rect 1400 2932 1452 2941
rect 7104 3136 7156 3188
rect 7288 3136 7340 3188
rect 3792 3111 3844 3120
rect 3792 3077 3801 3111
rect 3801 3077 3835 3111
rect 3835 3077 3844 3111
rect 3792 3068 3844 3077
rect 5632 3111 5684 3120
rect 5632 3077 5641 3111
rect 5641 3077 5675 3111
rect 5675 3077 5684 3111
rect 5632 3068 5684 3077
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 3148 3000 3200 3052
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3976 3043 4028 3052
rect 3700 3000 3752 3009
rect 3976 3009 3985 3043
rect 3985 3009 4019 3043
rect 4019 3009 4028 3043
rect 3976 3000 4028 3009
rect 4620 3043 4672 3052
rect 4620 3009 4629 3043
rect 4629 3009 4663 3043
rect 4663 3009 4672 3043
rect 4620 3000 4672 3009
rect 5080 3000 5132 3052
rect 5540 3043 5592 3052
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 5724 3000 5776 3052
rect 7656 3068 7708 3120
rect 8668 3136 8720 3188
rect 9220 3179 9272 3188
rect 9220 3145 9229 3179
rect 9229 3145 9263 3179
rect 9263 3145 9272 3179
rect 9220 3136 9272 3145
rect 9772 3136 9824 3188
rect 11152 3136 11204 3188
rect 11520 3136 11572 3188
rect 6828 2932 6880 2984
rect 1860 2864 1912 2916
rect 3792 2864 3844 2916
rect 5172 2864 5224 2916
rect 2780 2796 2832 2848
rect 4344 2796 4396 2848
rect 4804 2796 4856 2848
rect 5540 2864 5592 2916
rect 7104 2864 7156 2916
rect 7472 3000 7524 3052
rect 9036 3000 9088 3052
rect 11796 3068 11848 3120
rect 11060 3000 11112 3052
rect 11888 3000 11940 3052
rect 7932 2932 7984 2984
rect 9864 2975 9916 2984
rect 8944 2864 8996 2916
rect 9864 2941 9873 2975
rect 9873 2941 9907 2975
rect 9907 2941 9916 2975
rect 9864 2932 9916 2941
rect 11980 2932 12032 2984
rect 12900 3000 12952 3052
rect 13636 3043 13688 3052
rect 13636 3009 13645 3043
rect 13645 3009 13679 3043
rect 13679 3009 13688 3043
rect 13636 3000 13688 3009
rect 14648 2975 14700 2984
rect 14648 2941 14657 2975
rect 14657 2941 14691 2975
rect 14691 2941 14700 2975
rect 14648 2932 14700 2941
rect 9956 2864 10008 2916
rect 11152 2864 11204 2916
rect 12256 2864 12308 2916
rect 6736 2796 6788 2848
rect 7380 2796 7432 2848
rect 7932 2839 7984 2848
rect 7932 2805 7941 2839
rect 7941 2805 7975 2839
rect 7975 2805 7984 2839
rect 7932 2796 7984 2805
rect 9128 2796 9180 2848
rect 9496 2796 9548 2848
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 12072 2796 12124 2848
rect 12164 2796 12216 2848
rect 3420 2694 3472 2746
rect 3484 2694 3536 2746
rect 3548 2694 3600 2746
rect 3612 2694 3664 2746
rect 8296 2694 8348 2746
rect 8360 2694 8412 2746
rect 8424 2694 8476 2746
rect 8488 2694 8540 2746
rect 13172 2694 13224 2746
rect 13236 2694 13288 2746
rect 13300 2694 13352 2746
rect 13364 2694 13416 2746
rect 3148 2635 3200 2644
rect 3148 2601 3157 2635
rect 3157 2601 3191 2635
rect 3191 2601 3200 2635
rect 3148 2592 3200 2601
rect 4620 2592 4672 2644
rect 7196 2592 7248 2644
rect 2872 2524 2924 2576
rect 6920 2524 6972 2576
rect 9036 2524 9088 2576
rect 3056 2456 3108 2508
rect 4344 2499 4396 2508
rect 4344 2465 4353 2499
rect 4353 2465 4387 2499
rect 4387 2465 4396 2499
rect 4344 2456 4396 2465
rect 7196 2499 7248 2508
rect 20 2388 72 2440
rect 2780 2388 2832 2440
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 3240 2431 3292 2440
rect 2964 2388 3016 2397
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 4988 2320 5040 2372
rect 7196 2465 7205 2499
rect 7205 2465 7239 2499
rect 7239 2465 7248 2499
rect 7196 2456 7248 2465
rect 8024 2456 8076 2508
rect 11152 2592 11204 2644
rect 11244 2592 11296 2644
rect 12532 2592 12584 2644
rect 14648 2592 14700 2644
rect 9588 2524 9640 2576
rect 9864 2524 9916 2576
rect 7012 2431 7064 2440
rect 7012 2397 7021 2431
rect 7021 2397 7055 2431
rect 7055 2397 7064 2431
rect 7012 2388 7064 2397
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 13728 2524 13780 2576
rect 14372 2524 14424 2576
rect 14832 2524 14884 2576
rect 14924 2456 14976 2508
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9404 2431 9456 2440
rect 9036 2320 9088 2372
rect 9404 2397 9413 2431
rect 9413 2397 9447 2431
rect 9447 2397 9456 2431
rect 9404 2388 9456 2397
rect 11520 2431 11572 2440
rect 9312 2320 9364 2372
rect 10232 2363 10284 2372
rect 10232 2329 10241 2363
rect 10241 2329 10275 2363
rect 10275 2329 10284 2363
rect 10232 2320 10284 2329
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 11796 2431 11848 2440
rect 11796 2397 11805 2431
rect 11805 2397 11839 2431
rect 11839 2397 11848 2431
rect 11796 2388 11848 2397
rect 11980 2388 12032 2440
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 14740 2431 14792 2440
rect 13912 2320 13964 2372
rect 14372 2363 14424 2372
rect 14372 2329 14381 2363
rect 14381 2329 14415 2363
rect 14415 2329 14424 2363
rect 14372 2320 14424 2329
rect 14740 2397 14749 2431
rect 14749 2397 14783 2431
rect 14783 2397 14792 2431
rect 14740 2388 14792 2397
rect 14832 2431 14884 2440
rect 14832 2397 14841 2431
rect 14841 2397 14875 2431
rect 14875 2397 14884 2431
rect 14832 2388 14884 2397
rect 6828 2295 6880 2304
rect 6828 2261 6837 2295
rect 6837 2261 6871 2295
rect 6871 2261 6880 2295
rect 6828 2252 6880 2261
rect 7656 2252 7708 2304
rect 9220 2252 9272 2304
rect 16764 2320 16816 2372
rect 14740 2252 14792 2304
rect 5858 2150 5910 2202
rect 5922 2150 5974 2202
rect 5986 2150 6038 2202
rect 6050 2150 6102 2202
rect 10734 2150 10786 2202
rect 10798 2150 10850 2202
rect 10862 2150 10914 2202
rect 10926 2150 10978 2202
rect 6644 2048 6696 2100
rect 10232 2048 10284 2100
rect 10600 1912 10652 1964
rect 12900 1912 12952 1964
rect 10508 1096 10560 1148
rect 11060 1096 11112 1148
<< metal2 >>
rect 18 18215 74 19015
rect 1858 18215 1914 19015
rect 3882 18215 3938 19015
rect 5722 18215 5778 19015
rect 7562 18215 7618 19015
rect 9402 18215 9458 19015
rect 11242 18215 11298 19015
rect 13082 18215 13138 19015
rect 14922 18215 14978 19015
rect 16762 18215 16818 19015
rect 32 14890 60 18215
rect 1872 16574 1900 18215
rect 1872 16546 1992 16574
rect 1398 16416 1454 16425
rect 1398 16351 1454 16360
rect 1412 16114 1440 16351
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1596 15026 1624 15506
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1688 15026 1716 15438
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1872 15094 1900 15302
rect 1964 15162 1992 16546
rect 3896 16182 3924 18215
rect 3884 16176 3936 16182
rect 3884 16118 3936 16124
rect 5736 16114 5764 18215
rect 5832 16348 6128 16368
rect 5888 16346 5912 16348
rect 5968 16346 5992 16348
rect 6048 16346 6072 16348
rect 5910 16294 5912 16346
rect 5974 16294 5986 16346
rect 6048 16294 6050 16346
rect 5888 16292 5912 16294
rect 5968 16292 5992 16294
rect 6048 16292 6072 16294
rect 5832 16272 6128 16292
rect 7576 16182 7604 18215
rect 9416 16674 9444 18215
rect 9416 16646 9628 16674
rect 9600 16266 9628 16646
rect 10708 16348 11004 16368
rect 10764 16346 10788 16348
rect 10844 16346 10868 16348
rect 10924 16346 10948 16348
rect 10786 16294 10788 16346
rect 10850 16294 10862 16346
rect 10924 16294 10926 16346
rect 10764 16292 10788 16294
rect 10844 16292 10868 16294
rect 10924 16292 10948 16294
rect 10708 16272 11004 16292
rect 9600 16238 9720 16266
rect 9692 16182 9720 16238
rect 7564 16176 7616 16182
rect 7564 16118 7616 16124
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 11256 16114 11284 18215
rect 13096 16182 13124 18215
rect 13084 16176 13136 16182
rect 13084 16118 13136 16124
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2056 15570 2084 15846
rect 2884 15638 2912 16050
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 2976 15502 3004 16050
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 1860 15088 1912 15094
rect 1860 15030 1912 15036
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 20 14884 72 14890
rect 20 14826 72 14832
rect 1584 14816 1636 14822
rect 1584 14758 1636 14764
rect 1596 10826 1624 14758
rect 1688 14618 1716 14962
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 2056 14482 2084 14962
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 2240 14346 2268 14758
rect 2228 14340 2280 14346
rect 2228 14282 2280 14288
rect 2688 14340 2740 14346
rect 2688 14282 2740 14288
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1872 13705 1900 13874
rect 1858 13696 1914 13705
rect 1858 13631 1914 13640
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1688 12782 1716 13330
rect 2240 13138 2268 14282
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2424 13326 2452 13874
rect 2700 13530 2728 14282
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2240 13110 2360 13138
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 11898 1716 12718
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1964 11354 1992 11698
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 1858 10976 1914 10985
rect 1858 10911 1914 10920
rect 1596 10798 1716 10826
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1596 6798 1624 7686
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 6254 1624 6598
rect 1688 6458 1716 10798
rect 1872 10266 1900 10911
rect 2056 10810 2084 11154
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 2240 9994 2268 10610
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2332 9178 2360 13110
rect 2424 12986 2452 13262
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2792 12782 2820 13194
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2792 12442 2820 12718
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2504 10668 2556 10674
rect 2556 10628 2636 10656
rect 2504 10610 2556 10616
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2424 9518 2452 10542
rect 2608 9994 2636 10628
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2700 10130 2728 10406
rect 2884 10198 2912 15302
rect 3160 15026 3188 15846
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3160 14074 3188 14962
rect 3252 14958 3280 16050
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 3394 15804 3690 15824
rect 3450 15802 3474 15804
rect 3530 15802 3554 15804
rect 3610 15802 3634 15804
rect 3472 15750 3474 15802
rect 3536 15750 3548 15802
rect 3610 15750 3612 15802
rect 3450 15748 3474 15750
rect 3530 15748 3554 15750
rect 3610 15748 3634 15750
rect 3394 15728 3690 15748
rect 3424 15360 3476 15366
rect 3424 15302 3476 15308
rect 3436 15162 3464 15302
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3394 14716 3690 14736
rect 3450 14714 3474 14716
rect 3530 14714 3554 14716
rect 3610 14714 3634 14716
rect 3472 14662 3474 14714
rect 3536 14662 3548 14714
rect 3610 14662 3612 14714
rect 3450 14660 3474 14662
rect 3530 14660 3554 14662
rect 3610 14660 3634 14662
rect 3394 14640 3690 14660
rect 4080 14618 4108 14894
rect 4172 14890 4200 15914
rect 4160 14884 4212 14890
rect 4160 14826 4212 14832
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 3160 13326 3188 13806
rect 3394 13628 3690 13648
rect 3450 13626 3474 13628
rect 3530 13626 3554 13628
rect 3610 13626 3634 13628
rect 3472 13574 3474 13626
rect 3536 13574 3548 13626
rect 3610 13574 3612 13626
rect 3450 13572 3474 13574
rect 3530 13572 3554 13574
rect 3610 13572 3634 13574
rect 3394 13552 3690 13572
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3068 12238 3096 12786
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2976 11150 3004 11630
rect 3056 11620 3108 11626
rect 3056 11562 3108 11568
rect 3068 11354 3096 11562
rect 3160 11354 3188 13262
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 3394 12540 3690 12560
rect 3450 12538 3474 12540
rect 3530 12538 3554 12540
rect 3610 12538 3634 12540
rect 3472 12486 3474 12538
rect 3536 12486 3548 12538
rect 3610 12486 3612 12538
rect 3450 12484 3474 12486
rect 3530 12484 3554 12486
rect 3610 12484 3634 12486
rect 3394 12464 3690 12484
rect 4080 12238 4108 12582
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2608 9722 2636 9930
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2700 9654 2728 10066
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2976 9450 3004 11086
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 8294 1900 8842
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1872 7886 1900 8230
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 2148 7750 2176 8910
rect 3160 8566 3188 11018
rect 3252 10674 3280 11698
rect 3394 11452 3690 11472
rect 3450 11450 3474 11452
rect 3530 11450 3554 11452
rect 3610 11450 3634 11452
rect 3472 11398 3474 11450
rect 3536 11398 3548 11450
rect 3610 11398 3612 11450
rect 3450 11396 3474 11398
rect 3530 11396 3554 11398
rect 3610 11396 3634 11398
rect 3394 11376 3690 11396
rect 3804 11150 3832 11698
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3620 10810 3648 11086
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3394 10364 3690 10384
rect 3450 10362 3474 10364
rect 3530 10362 3554 10364
rect 3610 10362 3634 10364
rect 3472 10310 3474 10362
rect 3536 10310 3548 10362
rect 3610 10310 3612 10362
rect 3450 10308 3474 10310
rect 3530 10308 3554 10310
rect 3610 10308 3634 10310
rect 3394 10288 3690 10308
rect 3790 9480 3846 9489
rect 3790 9415 3846 9424
rect 3394 9276 3690 9296
rect 3450 9274 3474 9276
rect 3530 9274 3554 9276
rect 3610 9274 3634 9276
rect 3472 9222 3474 9274
rect 3536 9222 3548 9274
rect 3610 9222 3612 9274
rect 3450 9220 3474 9222
rect 3530 9220 3554 9222
rect 3610 9220 3634 9222
rect 3394 9200 3690 9220
rect 3804 8974 3832 9415
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 3896 8498 3924 11494
rect 3988 10266 4016 12174
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 4172 11150 4200 11698
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9722 4200 9998
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3988 8838 4016 8978
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2332 8090 2360 8366
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2688 7880 2740 7886
rect 2792 7868 2820 8434
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2884 8265 2912 8298
rect 3148 8288 3200 8294
rect 2870 8256 2926 8265
rect 3148 8230 3200 8236
rect 2870 8191 2926 8200
rect 3160 7954 3188 8230
rect 3394 8188 3690 8208
rect 3450 8186 3474 8188
rect 3530 8186 3554 8188
rect 3610 8186 3634 8188
rect 3472 8134 3474 8186
rect 3536 8134 3548 8186
rect 3610 8134 3612 8186
rect 3450 8132 3474 8134
rect 3530 8132 3554 8134
rect 3610 8132 3634 8134
rect 3394 8112 3690 8132
rect 3700 8016 3752 8022
rect 3700 7958 3752 7964
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 2740 7840 2820 7868
rect 2688 7822 2740 7828
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 3160 7478 3188 7890
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3712 7410 3740 7958
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 2884 7002 2912 7346
rect 3896 7342 3924 8434
rect 3988 7886 4016 8774
rect 4080 8566 4108 8774
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 4080 7410 4108 8502
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1596 5710 1624 6190
rect 1688 5710 1716 6394
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 2056 5914 2084 6054
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 2148 5710 2176 6802
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2332 5642 2360 6598
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2412 5704 2464 5710
rect 2410 5672 2412 5681
rect 2464 5672 2466 5681
rect 2320 5636 2372 5642
rect 2410 5607 2466 5616
rect 2320 5578 2372 5584
rect 2608 5574 2636 6122
rect 1584 5568 1636 5574
rect 1398 5536 1454 5545
rect 1584 5510 1636 5516
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 1398 5471 1454 5480
rect 1412 5234 1440 5471
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1596 4622 1624 5510
rect 2884 5370 2912 6938
rect 3252 6730 3280 7142
rect 3394 7100 3690 7120
rect 3450 7098 3474 7100
rect 3530 7098 3554 7100
rect 3610 7098 3634 7100
rect 3472 7046 3474 7098
rect 3536 7046 3548 7098
rect 3610 7046 3612 7098
rect 3450 7044 3474 7046
rect 3530 7044 3554 7046
rect 3610 7044 3634 7046
rect 3394 7024 3690 7044
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2424 5137 2452 5170
rect 2410 5128 2466 5137
rect 2410 5063 2466 5072
rect 2044 4752 2096 4758
rect 2044 4694 2096 4700
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 2056 4146 2084 4694
rect 3068 4622 3096 6598
rect 3252 6390 3280 6666
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 3252 5846 3280 6122
rect 3394 6012 3690 6032
rect 3450 6010 3474 6012
rect 3530 6010 3554 6012
rect 3610 6010 3634 6012
rect 3472 5958 3474 6010
rect 3536 5958 3548 6010
rect 3610 5958 3612 6010
rect 3450 5956 3474 5958
rect 3530 5956 3554 5958
rect 3610 5956 3634 5958
rect 3394 5936 3690 5956
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 3988 5778 4016 6734
rect 4080 6458 4108 6734
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4080 5710 4108 6394
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 3160 5234 3188 5306
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3976 5228 4028 5234
rect 4264 5216 4292 16050
rect 5080 14544 5132 14550
rect 5080 14486 5132 14492
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4724 13258 4752 14350
rect 4816 14074 4844 14350
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4816 13394 4844 14010
rect 4908 14006 4936 14214
rect 4896 14000 4948 14006
rect 4896 13942 4948 13948
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4712 13252 4764 13258
rect 4712 13194 4764 13200
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4356 12238 4384 12650
rect 4448 12306 4476 12718
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4448 10198 4476 12242
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4540 10674 4568 10950
rect 4908 10810 4936 13942
rect 5092 13938 5120 14486
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5092 12986 5120 13874
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5276 12434 5304 16050
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5460 15638 5488 15846
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5368 15162 5396 15302
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5460 14958 5488 15574
rect 5632 15428 5684 15434
rect 5632 15370 5684 15376
rect 6184 15428 6236 15434
rect 6184 15370 6236 15376
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 13870 5580 14350
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5644 13530 5672 15370
rect 5832 15260 6128 15280
rect 5888 15258 5912 15260
rect 5968 15258 5992 15260
rect 6048 15258 6072 15260
rect 5910 15206 5912 15258
rect 5974 15206 5986 15258
rect 6048 15206 6050 15258
rect 5888 15204 5912 15206
rect 5968 15204 5992 15206
rect 6048 15204 6072 15206
rect 5832 15184 6128 15204
rect 6196 15162 6224 15370
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 5832 14172 6128 14192
rect 5888 14170 5912 14172
rect 5968 14170 5992 14172
rect 6048 14170 6072 14172
rect 5910 14118 5912 14170
rect 5974 14118 5986 14170
rect 6048 14118 6050 14170
rect 5888 14116 5912 14118
rect 5968 14116 5992 14118
rect 6048 14116 6072 14118
rect 5832 14096 6128 14116
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5368 12442 5396 13262
rect 5736 12986 5764 13874
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 5828 13462 5856 13806
rect 6184 13796 6236 13802
rect 6184 13738 6236 13744
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5832 13084 6128 13104
rect 5888 13082 5912 13084
rect 5968 13082 5992 13084
rect 6048 13082 6072 13084
rect 5910 13030 5912 13082
rect 5974 13030 5986 13082
rect 6048 13030 6050 13082
rect 5888 13028 5912 13030
rect 5968 13028 5992 13030
rect 6048 13028 6072 13030
rect 5832 13008 6128 13028
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 6196 12850 6224 13738
rect 6564 12850 6592 15982
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 5092 12406 5304 12434
rect 5356 12436 5408 12442
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 5000 10810 5028 11018
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4632 9926 4660 10474
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4448 8974 4476 9454
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4448 6458 4476 6802
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4632 5302 4660 9862
rect 4908 9674 4936 9998
rect 4908 9654 5028 9674
rect 4908 9648 5040 9654
rect 4908 9646 4988 9648
rect 4988 9590 5040 9596
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4724 8974 4752 9386
rect 5000 8974 5028 9590
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4908 5234 4936 6326
rect 5000 6254 5028 6598
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5000 5234 5028 6190
rect 3976 5170 4028 5176
rect 4172 5188 4292 5216
rect 4344 5228 4396 5234
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 2136 4548 2188 4554
rect 2136 4490 2188 4496
rect 2148 4146 2176 4490
rect 2424 4146 2452 4558
rect 2964 4480 3016 4486
rect 3160 4434 3188 5170
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3394 4924 3690 4944
rect 3450 4922 3474 4924
rect 3530 4922 3554 4924
rect 3610 4922 3634 4924
rect 3472 4870 3474 4922
rect 3536 4870 3548 4922
rect 3610 4870 3612 4922
rect 3450 4868 3474 4870
rect 3530 4868 3554 4870
rect 3610 4868 3634 4870
rect 3394 4848 3690 4868
rect 2964 4422 3016 4428
rect 2976 4282 3004 4422
rect 3068 4406 3188 4434
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2976 4078 3004 4218
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1412 2825 1440 2926
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1398 2816 1454 2825
rect 1398 2751 1454 2760
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 32 800 60 2382
rect 1872 800 1900 2858
rect 2792 2854 2820 3538
rect 2976 3398 3004 3878
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2792 2446 2820 2790
rect 2884 2582 2912 2994
rect 2872 2576 2924 2582
rect 2872 2518 2924 2524
rect 2976 2446 3004 3334
rect 3068 2514 3096 4406
rect 3394 3836 3690 3856
rect 3450 3834 3474 3836
rect 3530 3834 3554 3836
rect 3610 3834 3634 3836
rect 3472 3782 3474 3834
rect 3536 3782 3548 3834
rect 3610 3782 3612 3834
rect 3450 3780 3474 3782
rect 3530 3780 3554 3782
rect 3610 3780 3634 3782
rect 3394 3760 3690 3780
rect 3804 3618 3832 4966
rect 3988 4826 4016 5170
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3988 4146 4016 4762
rect 4080 4758 4108 5034
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 4172 4690 4200 5188
rect 4344 5170 4396 5176
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4264 4570 4292 5034
rect 4356 4690 4384 5170
rect 4712 5024 4764 5030
rect 5092 5012 5120 12406
rect 5356 12378 5408 12384
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5644 11762 5672 12174
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5276 11354 5304 11698
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 10826 5580 11018
rect 5368 10798 5580 10826
rect 5368 10742 5396 10798
rect 5356 10736 5408 10742
rect 5356 10678 5408 10684
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5460 9178 5488 9454
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5460 8634 5488 9114
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5552 8514 5580 10678
rect 5644 10062 5672 11222
rect 5736 11150 5764 12786
rect 6564 12730 6592 12786
rect 6380 12702 6592 12730
rect 6380 12434 6408 12702
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6288 12406 6408 12434
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 5832 11996 6128 12016
rect 5888 11994 5912 11996
rect 5968 11994 5992 11996
rect 6048 11994 6072 11996
rect 5910 11942 5912 11994
rect 5974 11942 5986 11994
rect 6048 11942 6050 11994
rect 5888 11940 5912 11942
rect 5968 11940 5992 11942
rect 6048 11940 6072 11942
rect 5832 11920 6128 11940
rect 6196 11762 6224 12106
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 6288 11082 6316 12406
rect 6564 12238 6592 12582
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6564 11694 6592 12174
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6472 11354 6500 11630
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 5832 10908 6128 10928
rect 5888 10906 5912 10908
rect 5968 10906 5992 10908
rect 6048 10906 6072 10908
rect 5910 10854 5912 10906
rect 5974 10854 5986 10906
rect 6048 10854 6050 10906
rect 5888 10852 5912 10854
rect 5968 10852 5992 10854
rect 6048 10852 6072 10854
rect 5832 10832 6128 10852
rect 5722 10704 5778 10713
rect 5722 10639 5724 10648
rect 5776 10639 5778 10648
rect 5724 10610 5776 10616
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5832 9820 6128 9840
rect 5888 9818 5912 9820
rect 5968 9818 5992 9820
rect 6048 9818 6072 9820
rect 5910 9766 5912 9818
rect 5974 9766 5986 9818
rect 6048 9766 6050 9818
rect 5888 9764 5912 9766
rect 5968 9764 5992 9766
rect 6048 9764 6072 9766
rect 5832 9744 6128 9764
rect 5630 9616 5686 9625
rect 6288 9602 6316 11018
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6564 10112 6592 10746
rect 6380 10084 6592 10112
rect 6380 9722 6408 10084
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 5630 9551 5632 9560
rect 5684 9551 5686 9560
rect 5724 9580 5776 9586
rect 5632 9522 5684 9528
rect 6288 9574 6500 9602
rect 5724 9522 5776 9528
rect 5736 9489 5764 9522
rect 5722 9480 5778 9489
rect 5722 9415 5778 9424
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6380 9178 6408 9318
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 5832 8732 6128 8752
rect 5888 8730 5912 8732
rect 5968 8730 5992 8732
rect 6048 8730 6072 8732
rect 5910 8678 5912 8730
rect 5974 8678 5986 8730
rect 6048 8678 6050 8730
rect 5888 8676 5912 8678
rect 5968 8676 5992 8678
rect 6048 8676 6072 8678
rect 5832 8656 6128 8676
rect 5552 8486 5672 8514
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7954 5212 8230
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5184 7478 5212 7890
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5172 7472 5224 7478
rect 5172 7414 5224 7420
rect 5552 7342 5580 7754
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5276 6866 5304 7142
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5184 5166 5212 6734
rect 5276 5234 5304 6802
rect 5644 6322 5672 8486
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5736 8022 5764 8366
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5724 8016 5776 8022
rect 5724 7958 5776 7964
rect 5736 7206 5764 7958
rect 5920 7818 5948 8298
rect 5908 7812 5960 7818
rect 6276 7812 6328 7818
rect 5908 7754 5960 7760
rect 6196 7772 6276 7800
rect 5832 7644 6128 7664
rect 5888 7642 5912 7644
rect 5968 7642 5992 7644
rect 6048 7642 6072 7644
rect 5910 7590 5912 7642
rect 5974 7590 5986 7642
rect 6048 7590 6050 7642
rect 5888 7588 5912 7590
rect 5968 7588 5992 7590
rect 6048 7588 6072 7590
rect 5832 7568 6128 7588
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5832 6556 6128 6576
rect 5888 6554 5912 6556
rect 5968 6554 5992 6556
rect 6048 6554 6072 6556
rect 5910 6502 5912 6554
rect 5974 6502 5986 6554
rect 6048 6502 6050 6554
rect 5888 6500 5912 6502
rect 5968 6500 5992 6502
rect 6048 6500 6072 6502
rect 5832 6480 6128 6500
rect 5632 6316 5684 6322
rect 5684 6276 5764 6304
rect 5632 6258 5684 6264
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5092 4984 5212 5012
rect 4712 4966 4764 4972
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4724 4622 4752 4966
rect 4712 4616 4764 4622
rect 4264 4542 4384 4570
rect 4712 4558 4764 4564
rect 4356 4486 4384 4542
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4214 4384 4422
rect 4724 4282 4752 4558
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5092 3670 5120 3878
rect 3712 3590 3832 3618
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 4988 3596 5040 3602
rect 3712 3534 3740 3590
rect 4988 3538 5040 3544
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3160 2650 3188 2994
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3252 2446 3280 3470
rect 3608 3460 3660 3466
rect 3608 3402 3660 3408
rect 3620 3058 3648 3402
rect 3712 3058 3740 3470
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3804 3126 3832 3334
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3988 3058 4016 3470
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 3792 2916 3844 2922
rect 3792 2858 3844 2864
rect 3394 2748 3690 2768
rect 3450 2746 3474 2748
rect 3530 2746 3554 2748
rect 3610 2746 3634 2748
rect 3472 2694 3474 2746
rect 3536 2694 3548 2746
rect 3610 2694 3612 2746
rect 3450 2692 3474 2694
rect 3530 2692 3554 2694
rect 3610 2692 3634 2694
rect 3394 2672 3690 2692
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3804 1442 3832 2858
rect 4172 2446 4200 3402
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4356 2514 4384 2790
rect 4632 2650 4660 2994
rect 4816 2854 4844 3470
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4344 2508 4396 2514
rect 4344 2450 4396 2456
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 5000 2378 5028 3538
rect 5092 3058 5120 3606
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5184 2922 5212 4984
rect 5368 3534 5396 5646
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5368 3040 5396 3470
rect 5644 3126 5672 5510
rect 5736 4622 5764 6276
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6012 5710 6040 6054
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 5832 5468 6128 5488
rect 5888 5466 5912 5468
rect 5968 5466 5992 5468
rect 6048 5466 6072 5468
rect 5910 5414 5912 5466
rect 5974 5414 5986 5466
rect 6048 5414 6050 5466
rect 5888 5412 5912 5414
rect 5968 5412 5992 5414
rect 6048 5412 6072 5414
rect 5832 5392 6128 5412
rect 6196 5273 6224 7772
rect 6276 7754 6328 7760
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 6322 6316 6734
rect 6380 6390 6408 8434
rect 6472 7818 6500 9574
rect 6564 8906 6592 9930
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6380 6186 6408 6326
rect 6368 6180 6420 6186
rect 6368 6122 6420 6128
rect 6182 5264 6238 5273
rect 6182 5199 6238 5208
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5832 4380 6128 4400
rect 5888 4378 5912 4380
rect 5968 4378 5992 4380
rect 6048 4378 6072 4380
rect 5910 4326 5912 4378
rect 5974 4326 5986 4378
rect 6048 4326 6050 4378
rect 5888 4324 5912 4326
rect 5968 4324 5992 4326
rect 6048 4324 6072 4326
rect 5832 4304 6128 4324
rect 6196 4214 6224 5199
rect 6564 5166 6592 8842
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6288 4457 6316 4694
rect 6564 4622 6592 5102
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6274 4448 6330 4457
rect 6274 4383 6330 4392
rect 6380 4282 6408 4558
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6184 4208 6236 4214
rect 6184 4150 6236 4156
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5736 3058 5764 3946
rect 6380 3534 6408 4218
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6472 3534 6500 3606
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5832 3292 6128 3312
rect 5888 3290 5912 3292
rect 5968 3290 5992 3292
rect 6048 3290 6072 3292
rect 5910 3238 5912 3290
rect 5974 3238 5986 3290
rect 6048 3238 6050 3290
rect 5888 3236 5912 3238
rect 5968 3236 5992 3238
rect 6048 3236 6072 3238
rect 5832 3216 6128 3236
rect 5540 3052 5592 3058
rect 5368 3012 5540 3040
rect 5540 2994 5592 3000
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5172 2916 5224 2922
rect 5172 2858 5224 2864
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 3712 1414 3832 1442
rect 3712 800 3740 1414
rect 5552 800 5580 2858
rect 5832 2204 6128 2224
rect 5888 2202 5912 2204
rect 5968 2202 5992 2204
rect 6048 2202 6072 2204
rect 5910 2150 5912 2202
rect 5974 2150 5986 2202
rect 6048 2150 6050 2202
rect 5888 2148 5912 2150
rect 5968 2148 5992 2150
rect 6048 2148 6072 2150
rect 5832 2128 6128 2148
rect 6656 2106 6684 14758
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6748 11830 6776 13874
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6840 10810 6868 15982
rect 8270 15804 8566 15824
rect 8326 15802 8350 15804
rect 8406 15802 8430 15804
rect 8486 15802 8510 15804
rect 8348 15750 8350 15802
rect 8412 15750 8424 15802
rect 8486 15750 8488 15802
rect 8326 15748 8350 15750
rect 8406 15748 8430 15750
rect 8486 15748 8510 15750
rect 8270 15728 8566 15748
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7392 15026 7420 15438
rect 7944 15094 7972 15438
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7392 14618 7420 14962
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7576 14346 7604 14758
rect 7668 14550 7696 14962
rect 7944 14618 7972 15030
rect 9140 14958 9168 16050
rect 9232 15706 9260 16050
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9232 15162 9260 15642
rect 9416 15570 9444 15846
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9784 15434 9812 16050
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 10152 15162 10180 16050
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10324 15428 10376 15434
rect 10324 15370 10376 15376
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 8270 14716 8566 14736
rect 8326 14714 8350 14716
rect 8406 14714 8430 14716
rect 8486 14714 8510 14716
rect 8348 14662 8350 14714
rect 8412 14662 8424 14714
rect 8486 14662 8488 14714
rect 8326 14660 8350 14662
rect 8406 14660 8430 14662
rect 8486 14660 8510 14662
rect 8270 14640 8566 14660
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7024 12782 7052 13262
rect 7116 12850 7144 13670
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 7024 11898 7052 12718
rect 7208 12442 7236 13466
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7116 11778 7144 12242
rect 7024 11762 7144 11778
rect 7012 11756 7144 11762
rect 7064 11750 7144 11756
rect 7012 11698 7064 11704
rect 7024 11336 7052 11698
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7104 11348 7156 11354
rect 7024 11308 7104 11336
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6748 7886 6776 10474
rect 7024 9994 7052 11308
rect 7104 11290 7156 11296
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 8974 6960 9862
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7024 9178 7052 9522
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6932 8566 6960 8910
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6932 8072 6960 8502
rect 6932 8044 7052 8072
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 6730 6776 7822
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6840 6798 6868 7754
rect 6932 7546 6960 7890
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 7024 7410 7052 8044
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 7116 6497 7144 10950
rect 7208 10713 7236 11494
rect 7300 10962 7328 14214
rect 7576 14074 7604 14282
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8036 13530 8064 13806
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8024 12912 8076 12918
rect 8024 12854 8076 12860
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7484 12238 7512 12786
rect 8036 12442 8064 12854
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7392 12102 7420 12174
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7392 11762 7420 12038
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7392 11218 7420 11698
rect 7484 11286 7512 12174
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7300 10934 7420 10962
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7194 10704 7250 10713
rect 7194 10639 7196 10648
rect 7248 10639 7250 10648
rect 7196 10610 7248 10616
rect 7208 10579 7236 10610
rect 7300 9994 7328 10746
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7392 9674 7420 10934
rect 7484 10606 7512 11018
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7208 9646 7420 9674
rect 7102 6488 7158 6497
rect 7102 6423 7158 6432
rect 7116 6390 7144 6423
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 7104 6384 7156 6390
rect 7208 6361 7236 9646
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7300 8974 7328 9454
rect 7484 9042 7512 10542
rect 7576 10538 7604 11018
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7392 8922 7420 8978
rect 7392 8894 7512 8922
rect 7484 8838 7512 8894
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7392 8294 7420 8774
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7576 7886 7604 10474
rect 7668 10062 7696 12378
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7760 10062 7788 11562
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7852 10674 7880 11086
rect 7944 11082 7972 11698
rect 8036 11558 8064 11834
rect 8128 11762 8156 14214
rect 9312 14000 9364 14006
rect 9416 13988 9444 14214
rect 9364 13960 9444 13988
rect 9312 13942 9364 13948
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8270 13628 8566 13648
rect 8326 13626 8350 13628
rect 8406 13626 8430 13628
rect 8486 13626 8510 13628
rect 8348 13574 8350 13626
rect 8412 13574 8424 13626
rect 8486 13574 8488 13626
rect 8326 13572 8350 13574
rect 8406 13572 8430 13574
rect 8486 13572 8510 13574
rect 8270 13552 8566 13572
rect 8956 13530 8984 13874
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 8956 13258 8984 13466
rect 9220 13320 9272 13326
rect 9140 13280 9220 13308
rect 8944 13252 8996 13258
rect 8944 13194 8996 13200
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8270 12540 8566 12560
rect 8326 12538 8350 12540
rect 8406 12538 8430 12540
rect 8486 12538 8510 12540
rect 8348 12486 8350 12538
rect 8412 12486 8424 12538
rect 8486 12486 8488 12538
rect 8326 12484 8350 12486
rect 8406 12484 8430 12486
rect 8486 12484 8510 12486
rect 8270 12464 8566 12484
rect 8680 12442 8708 12650
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8668 12436 8720 12442
rect 8864 12434 8892 12582
rect 8668 12378 8720 12384
rect 8772 12406 8892 12434
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8312 12238 8340 12310
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8496 11898 8524 12242
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8270 11452 8566 11472
rect 8326 11450 8350 11452
rect 8406 11450 8430 11452
rect 8486 11450 8510 11452
rect 8348 11398 8350 11450
rect 8412 11398 8424 11450
rect 8486 11398 8488 11450
rect 8326 11396 8350 11398
rect 8406 11396 8430 11398
rect 8486 11396 8510 11398
rect 8270 11376 8566 11396
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7668 9586 7696 9998
rect 7760 9926 7788 9998
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7300 6866 7328 7278
rect 7484 7206 7512 7686
rect 7852 7478 7880 10610
rect 7932 10532 7984 10538
rect 7932 10474 7984 10480
rect 7944 10062 7972 10474
rect 8128 10470 8156 11222
rect 8680 11218 8708 12378
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8128 10062 8156 10406
rect 8270 10364 8566 10384
rect 8326 10362 8350 10364
rect 8406 10362 8430 10364
rect 8486 10362 8510 10364
rect 8348 10310 8350 10362
rect 8412 10310 8424 10362
rect 8486 10310 8488 10362
rect 8326 10308 8350 10310
rect 8406 10308 8430 10310
rect 8486 10308 8510 10310
rect 8270 10288 8566 10308
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7944 9586 7972 9998
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 8114 9480 8170 9489
rect 8114 9415 8170 9424
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7944 8974 7972 9318
rect 8128 9178 8156 9415
rect 8270 9276 8566 9296
rect 8326 9274 8350 9276
rect 8406 9274 8430 9276
rect 8486 9274 8510 9276
rect 8348 9222 8350 9274
rect 8412 9222 8424 9274
rect 8486 9222 8488 9274
rect 8326 9220 8350 9222
rect 8406 9220 8430 9222
rect 8486 9220 8510 9222
rect 8270 9200 8566 9220
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 8680 8498 8708 10406
rect 8772 9178 8800 12406
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9048 11694 9076 12174
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8864 10266 8892 11086
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8956 10674 8984 10950
rect 9048 10742 9076 11630
rect 9140 10810 9168 13280
rect 9220 13262 9272 13268
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9232 12442 9260 12786
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9324 12238 9352 13942
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9508 12782 9536 13874
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9508 12434 9536 12718
rect 9416 12406 9536 12434
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8956 8906 8984 10610
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 9048 9674 9076 9930
rect 9048 9646 9168 9674
rect 9140 9518 9168 9646
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8956 8498 8984 8842
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8270 8188 8566 8208
rect 8326 8186 8350 8188
rect 8406 8186 8430 8188
rect 8486 8186 8510 8188
rect 8348 8134 8350 8186
rect 8412 8134 8424 8186
rect 8486 8134 8488 8186
rect 8326 8132 8350 8134
rect 8406 8132 8430 8134
rect 8486 8132 8510 8134
rect 8270 8112 8566 8132
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7484 6882 7512 7142
rect 7576 6984 7604 7346
rect 7576 6956 7696 6984
rect 7288 6860 7340 6866
rect 7484 6854 7604 6882
rect 7668 6866 7696 6956
rect 7288 6802 7340 6808
rect 7576 6798 7604 6854
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7852 6798 7880 7414
rect 8270 7100 8566 7120
rect 8326 7098 8350 7100
rect 8406 7098 8430 7100
rect 8486 7098 8510 7100
rect 8348 7046 8350 7098
rect 8412 7046 8424 7098
rect 8486 7046 8488 7098
rect 8326 7044 8350 7046
rect 8406 7044 8430 7046
rect 8486 7044 8510 7046
rect 8270 7024 8566 7044
rect 8680 6798 8708 8434
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 7576 6662 7604 6734
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7104 6326 7156 6332
rect 7194 6352 7250 6361
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6748 2854 6776 5578
rect 6840 4593 6868 6326
rect 7194 6287 7196 6296
rect 7248 6287 7250 6296
rect 7196 6258 7248 6264
rect 7208 6227 7236 6258
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6932 5370 6960 5646
rect 7116 5642 7144 6054
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 7012 5228 7064 5234
rect 7116 5216 7144 5578
rect 7064 5188 7144 5216
rect 7012 5170 7064 5176
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6826 4584 6882 4593
rect 6826 4519 6882 4528
rect 7024 4146 7052 4626
rect 7392 4622 7420 5782
rect 7576 5098 7604 6598
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7852 4690 7880 5510
rect 7944 5216 7972 6734
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8036 5710 8064 6190
rect 8128 5710 8156 6326
rect 8404 6225 8432 6734
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8574 6624 8630 6633
rect 8496 6390 8524 6598
rect 8574 6559 8630 6568
rect 8588 6390 8616 6559
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 8390 6216 8446 6225
rect 8390 6151 8446 6160
rect 8270 6012 8566 6032
rect 8326 6010 8350 6012
rect 8406 6010 8430 6012
rect 8486 6010 8510 6012
rect 8348 5958 8350 6010
rect 8412 5958 8424 6010
rect 8486 5958 8488 6010
rect 8326 5956 8350 5958
rect 8406 5956 8430 5958
rect 8486 5956 8510 5958
rect 8270 5936 8566 5956
rect 8680 5760 8708 6734
rect 8496 5732 8708 5760
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8116 5704 8168 5710
rect 8392 5704 8444 5710
rect 8116 5646 8168 5652
rect 8206 5672 8262 5681
rect 8496 5692 8524 5732
rect 8444 5664 8524 5692
rect 8392 5646 8444 5652
rect 8206 5607 8262 5616
rect 8220 5574 8248 5607
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8772 5234 8800 8366
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8864 6458 8892 6938
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8956 6118 8984 7142
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8850 5264 8906 5273
rect 8024 5228 8076 5234
rect 7944 5188 8024 5216
rect 8024 5170 8076 5176
rect 8760 5228 8812 5234
rect 8956 5234 8984 6054
rect 8850 5199 8906 5208
rect 8944 5228 8996 5234
rect 8760 5170 8812 5176
rect 8036 4826 8064 5170
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 8128 4622 8156 5034
rect 8270 4924 8566 4944
rect 8326 4922 8350 4924
rect 8406 4922 8430 4924
rect 8486 4922 8510 4924
rect 8348 4870 8350 4922
rect 8412 4870 8424 4922
rect 8486 4870 8488 4922
rect 8326 4868 8350 4870
rect 8406 4868 8430 4870
rect 8486 4868 8510 4870
rect 8270 4848 8566 4868
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 8116 4616 8168 4622
rect 8680 4593 8708 4626
rect 8116 4558 8168 4564
rect 8666 4584 8722 4593
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7116 4146 7144 4422
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7392 4026 7420 4558
rect 8666 4519 8722 4528
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8220 4146 8248 4422
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 7300 4010 7420 4026
rect 7288 4004 7420 4010
rect 7340 3998 7420 4004
rect 7288 3946 7340 3952
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6840 2310 6868 2926
rect 6932 2582 6960 3538
rect 7484 3534 7512 3878
rect 8270 3836 8566 3856
rect 8326 3834 8350 3836
rect 8406 3834 8430 3836
rect 8486 3834 8510 3836
rect 8348 3782 8350 3834
rect 8412 3782 8424 3834
rect 8486 3782 8488 3834
rect 8326 3780 8350 3782
rect 8406 3780 8430 3782
rect 8486 3780 8510 3782
rect 8270 3760 8566 3780
rect 8680 3670 8708 4082
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7012 3528 7064 3534
rect 7010 3496 7012 3505
rect 7196 3528 7248 3534
rect 7064 3496 7066 3505
rect 7196 3470 7248 3476
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7010 3431 7066 3440
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 7024 2446 7052 3431
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7116 3194 7144 3334
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7102 2952 7158 2961
rect 7102 2887 7104 2896
rect 7156 2887 7158 2896
rect 7104 2858 7156 2864
rect 7208 2650 7236 3470
rect 7300 3194 7328 3470
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7484 3058 7512 3470
rect 7668 3466 7696 3538
rect 8116 3528 8168 3534
rect 8114 3496 8116 3505
rect 8168 3496 8170 3505
rect 7656 3460 7708 3466
rect 8114 3431 8170 3440
rect 7656 3402 7708 3408
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 7852 3074 7880 3334
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7208 2514 7236 2586
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 7392 800 7420 2790
rect 7668 2310 7696 3062
rect 7852 3046 7972 3074
rect 7944 2990 7972 3046
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 7944 2446 7972 2790
rect 8036 2514 8064 3334
rect 8680 3194 8708 3606
rect 8772 3534 8800 5170
rect 8864 4758 8892 5199
rect 8944 5170 8996 5176
rect 8956 5098 8984 5170
rect 8944 5092 8996 5098
rect 8944 5034 8996 5040
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 8944 4548 8996 4554
rect 8944 4490 8996 4496
rect 8956 4282 8984 4490
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 9048 4026 9076 9114
rect 9140 6186 9168 9454
rect 9232 8566 9260 11494
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9324 10062 9352 11018
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9324 9722 9352 9998
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9416 9489 9444 12406
rect 9600 10674 9628 14282
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9784 12374 9812 12786
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9876 12322 9904 14350
rect 10336 14074 10364 15370
rect 10428 14618 10456 15438
rect 10508 15428 10560 15434
rect 10508 15370 10560 15376
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10428 14006 10456 14554
rect 10416 14000 10468 14006
rect 10416 13942 10468 13948
rect 10520 13938 10548 15370
rect 10708 15260 11004 15280
rect 10764 15258 10788 15260
rect 10844 15258 10868 15260
rect 10924 15258 10948 15260
rect 10786 15206 10788 15258
rect 10850 15206 10862 15258
rect 10924 15206 10926 15258
rect 10764 15204 10788 15206
rect 10844 15204 10868 15206
rect 10924 15204 10948 15206
rect 10708 15184 11004 15204
rect 11060 14340 11112 14346
rect 11060 14282 11112 14288
rect 10708 14172 11004 14192
rect 10764 14170 10788 14172
rect 10844 14170 10868 14172
rect 10924 14170 10948 14172
rect 10786 14118 10788 14170
rect 10850 14118 10862 14170
rect 10924 14118 10926 14170
rect 10764 14116 10788 14118
rect 10844 14116 10868 14118
rect 10924 14116 10948 14118
rect 10708 14096 11004 14116
rect 11072 13988 11100 14282
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11164 14006 11192 14214
rect 10980 13960 11100 13988
rect 11152 14000 11204 14006
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10876 13932 10928 13938
rect 10980 13920 11008 13960
rect 11152 13942 11204 13948
rect 11716 13938 11744 15846
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11808 14414 11836 15302
rect 12084 14958 12112 15438
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12268 15026 12296 15370
rect 12636 15162 12664 15982
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12268 14618 12296 14962
rect 12820 14906 12848 15846
rect 13146 15804 13442 15824
rect 13202 15802 13226 15804
rect 13282 15802 13306 15804
rect 13362 15802 13386 15804
rect 13224 15750 13226 15802
rect 13288 15750 13300 15802
rect 13362 15750 13364 15802
rect 13202 15748 13226 15750
rect 13282 15748 13306 15750
rect 13362 15748 13386 15750
rect 13146 15728 13442 15748
rect 12900 15632 12952 15638
rect 12900 15574 12952 15580
rect 12912 15026 12940 15574
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12820 14878 12940 14906
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12440 14544 12492 14550
rect 12440 14486 12492 14492
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 11704 13932 11756 13938
rect 10928 13892 11008 13920
rect 11624 13892 11704 13920
rect 10876 13874 10928 13880
rect 10888 13326 10916 13874
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 10060 12918 10088 13194
rect 10048 12912 10100 12918
rect 10048 12854 10100 12860
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9968 12442 9996 12786
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 9876 12306 9996 12322
rect 9876 12300 10008 12306
rect 9876 12294 9956 12300
rect 9956 12242 10008 12248
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9784 11830 9812 12174
rect 9968 11898 9996 12242
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 10060 11234 10088 12854
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10152 12102 10180 12582
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10152 11898 10180 12038
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 9784 10742 9812 11222
rect 10060 11206 10180 11234
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9600 9874 9628 10610
rect 9680 10124 9732 10130
rect 9784 10112 9812 10678
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9732 10084 9812 10112
rect 9680 10066 9732 10072
rect 9876 10062 9904 10542
rect 10060 10266 10088 11018
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9600 9846 9720 9874
rect 9588 9716 9640 9722
rect 9508 9676 9588 9704
rect 9508 9518 9536 9676
rect 9588 9658 9640 9664
rect 9692 9602 9720 9846
rect 9600 9574 9720 9602
rect 9496 9512 9548 9518
rect 9402 9480 9458 9489
rect 9312 9444 9364 9450
rect 9496 9454 9548 9460
rect 9402 9415 9458 9424
rect 9312 9386 9364 9392
rect 9324 9178 9352 9386
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9416 9024 9444 9415
rect 9324 8996 9444 9024
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9324 8362 9352 8996
rect 9600 8922 9628 9574
rect 9680 9512 9732 9518
rect 9678 9480 9680 9489
rect 9732 9480 9734 9489
rect 9678 9415 9734 9424
rect 9416 8894 9628 8922
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 9140 6089 9168 6122
rect 9126 6080 9182 6089
rect 9126 6015 9182 6024
rect 9232 5914 9260 6734
rect 9416 6610 9444 8894
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9600 8498 9628 8774
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9508 7818 9536 8366
rect 9600 7886 9628 8434
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9692 7562 9720 9415
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9876 8362 9904 8910
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9600 7534 9720 7562
rect 9600 6633 9628 7534
rect 9876 7410 9904 8298
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9876 6798 9904 7346
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9413 6582 9444 6610
rect 9586 6624 9642 6633
rect 9413 6440 9441 6582
rect 9586 6559 9642 6568
rect 9586 6488 9642 6497
rect 9413 6412 9444 6440
rect 9586 6423 9588 6432
rect 9312 6384 9364 6390
rect 9310 6352 9312 6361
rect 9364 6352 9366 6361
rect 9310 6287 9366 6296
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9140 5030 9168 5170
rect 9324 5114 9352 6122
rect 9416 5234 9444 6412
rect 9640 6423 9642 6432
rect 9588 6394 9640 6400
rect 9968 6322 9996 8230
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10060 7546 10088 7754
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10152 7206 10180 11206
rect 10244 11082 10272 13262
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10336 11558 10364 13126
rect 10508 12912 10560 12918
rect 10428 12872 10508 12900
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 10428 10742 10456 12872
rect 10508 12854 10560 12860
rect 10612 11354 10640 13262
rect 10708 13084 11004 13104
rect 10764 13082 10788 13084
rect 10844 13082 10868 13084
rect 10924 13082 10948 13084
rect 10786 13030 10788 13082
rect 10850 13030 10862 13082
rect 10924 13030 10926 13082
rect 10764 13028 10788 13030
rect 10844 13028 10868 13030
rect 10924 13028 10948 13030
rect 10708 13008 11004 13028
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10704 12238 10732 12718
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10708 11996 11004 12016
rect 10764 11994 10788 11996
rect 10844 11994 10868 11996
rect 10924 11994 10948 11996
rect 10786 11942 10788 11994
rect 10850 11942 10862 11994
rect 10924 11942 10926 11994
rect 10764 11940 10788 11942
rect 10844 11940 10868 11942
rect 10924 11940 10948 11942
rect 10708 11920 11004 11940
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10704 11558 10732 11766
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10508 11076 10560 11082
rect 10704 11064 10732 11494
rect 10508 11018 10560 11024
rect 10612 11036 10732 11064
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10244 7410 10272 9862
rect 10428 9722 10456 10678
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10244 6730 10272 7346
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9588 6248 9640 6254
rect 9586 6216 9588 6225
rect 9640 6216 9642 6225
rect 9496 6180 9548 6186
rect 9586 6151 9642 6160
rect 10140 6180 10192 6186
rect 9496 6122 9548 6128
rect 10140 6122 10192 6128
rect 9508 6089 9536 6122
rect 9494 6080 9550 6089
rect 9494 6015 9550 6024
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 9770 5672 9826 5681
rect 9770 5607 9772 5616
rect 9824 5607 9826 5616
rect 9772 5578 9824 5584
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9232 5086 9352 5114
rect 9404 5092 9456 5098
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9232 4622 9260 5086
rect 9404 5034 9456 5040
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9220 4616 9272 4622
rect 9140 4576 9220 4604
rect 9140 4146 9168 4576
rect 9220 4558 9272 4564
rect 9324 4214 9352 4966
rect 9416 4486 9444 5034
rect 9692 4690 9720 5510
rect 9876 5370 9904 5782
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9784 5137 9812 5306
rect 10060 5234 10088 5782
rect 10152 5574 10180 6122
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10152 5234 10180 5510
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9770 5128 9826 5137
rect 9770 5063 9826 5072
rect 10152 4978 10180 5170
rect 9968 4950 10180 4978
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9220 4140 9272 4146
rect 9416 4128 9444 4422
rect 9600 4282 9628 4558
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9692 4457 9720 4490
rect 9678 4448 9734 4457
rect 9678 4383 9734 4392
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 9416 4100 9628 4128
rect 9220 4082 9272 4088
rect 8956 3998 9076 4026
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8956 2922 8984 3998
rect 9232 3194 9260 4082
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8944 2916 8996 2922
rect 8944 2858 8996 2864
rect 8270 2748 8566 2768
rect 8326 2746 8350 2748
rect 8406 2746 8430 2748
rect 8486 2746 8510 2748
rect 8348 2694 8350 2746
rect 8412 2694 8424 2746
rect 8486 2694 8488 2746
rect 8326 2692 8350 2694
rect 8406 2692 8430 2694
rect 8486 2692 8510 2694
rect 8270 2672 8566 2692
rect 9048 2582 9076 2994
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9036 2576 9088 2582
rect 9036 2518 9088 2524
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 9048 2378 9076 2518
rect 9140 2446 9168 2790
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9232 2394 9260 3130
rect 9416 2446 9444 3946
rect 9508 2854 9536 4100
rect 9600 4026 9628 4100
rect 9600 3998 9904 4026
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9600 3602 9628 3878
rect 9876 3602 9904 3998
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9600 2582 9628 3538
rect 9680 3528 9732 3534
rect 9732 3476 9812 3482
rect 9680 3470 9812 3476
rect 9692 3454 9812 3470
rect 9784 3194 9812 3454
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9784 2854 9812 3130
rect 9876 2990 9904 3402
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9876 2582 9904 2926
rect 9968 2922 9996 4950
rect 10244 4554 10272 6666
rect 10336 6186 10364 9522
rect 10428 8906 10456 9658
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10520 8634 10548 11018
rect 10612 10656 10640 11036
rect 10708 10908 11004 10928
rect 10764 10906 10788 10908
rect 10844 10906 10868 10908
rect 10924 10906 10948 10908
rect 10786 10854 10788 10906
rect 10850 10854 10862 10906
rect 10924 10854 10926 10906
rect 10764 10852 10788 10854
rect 10844 10852 10868 10854
rect 10924 10852 10948 10854
rect 10708 10832 11004 10852
rect 10692 10668 10744 10674
rect 10612 10628 10692 10656
rect 10612 10470 10640 10628
rect 10692 10610 10744 10616
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 11072 10062 11100 13670
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11164 11898 11192 12174
rect 11348 11898 11376 13262
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11164 11150 11192 11630
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10708 9820 11004 9840
rect 10764 9818 10788 9820
rect 10844 9818 10868 9820
rect 10924 9818 10948 9820
rect 10786 9766 10788 9818
rect 10850 9766 10862 9818
rect 10924 9766 10926 9818
rect 10764 9764 10788 9766
rect 10844 9764 10868 9766
rect 10924 9764 10948 9766
rect 10708 9744 11004 9764
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10508 8628 10560 8634
rect 10612 8616 10640 9454
rect 11072 9382 11100 9998
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11164 9625 11192 9658
rect 11150 9616 11206 9625
rect 11150 9551 11206 9560
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 10708 8732 11004 8752
rect 10764 8730 10788 8732
rect 10844 8730 10868 8732
rect 10924 8730 10948 8732
rect 10786 8678 10788 8730
rect 10850 8678 10862 8730
rect 10924 8678 10926 8730
rect 10764 8676 10788 8678
rect 10844 8676 10868 8678
rect 10924 8676 10948 8678
rect 10708 8656 11004 8676
rect 10612 8588 10732 8616
rect 10508 8570 10560 8576
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10428 8022 10456 8434
rect 10506 8120 10562 8129
rect 10612 8090 10640 8434
rect 10704 8294 10732 8588
rect 11072 8566 11100 9046
rect 11256 8634 11284 9862
rect 11440 9178 11468 12106
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11532 11218 11560 11698
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11532 10470 11560 11154
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10506 8055 10508 8064
rect 10560 8055 10562 8064
rect 10600 8084 10652 8090
rect 10508 8026 10560 8032
rect 10600 8026 10652 8032
rect 10416 8016 10468 8022
rect 10704 7970 10732 8230
rect 10416 7958 10468 7964
rect 10612 7942 10732 7970
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10428 7546 10456 7822
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10612 7002 10640 7942
rect 11072 7886 11100 8366
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 10708 7644 11004 7664
rect 10764 7642 10788 7644
rect 10844 7642 10868 7644
rect 10924 7642 10948 7644
rect 10786 7590 10788 7642
rect 10850 7590 10862 7642
rect 10924 7590 10926 7642
rect 10764 7588 10788 7590
rect 10844 7588 10868 7590
rect 10924 7588 10948 7590
rect 10708 7568 11004 7588
rect 11164 7410 11192 7822
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10980 7002 11008 7278
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11072 7002 11100 7142
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10336 5234 10364 5510
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10336 4826 10364 5170
rect 10428 5098 10456 6802
rect 10708 6556 11004 6576
rect 10764 6554 10788 6556
rect 10844 6554 10868 6556
rect 10924 6554 10948 6556
rect 10786 6502 10788 6554
rect 10850 6502 10862 6554
rect 10924 6502 10926 6554
rect 10764 6500 10788 6502
rect 10844 6500 10868 6502
rect 10924 6500 10948 6502
rect 10708 6480 11004 6500
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10796 5710 10824 6258
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10784 5704 10836 5710
rect 10888 5692 10916 6054
rect 10980 5817 11008 6054
rect 10966 5808 11022 5817
rect 10966 5743 11022 5752
rect 10968 5704 11020 5710
rect 10888 5664 10968 5692
rect 10784 5646 10836 5652
rect 10968 5646 11020 5652
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10520 5370 10548 5578
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10612 5166 10640 5646
rect 10708 5468 11004 5488
rect 10764 5466 10788 5468
rect 10844 5466 10868 5468
rect 10924 5466 10948 5468
rect 10786 5414 10788 5466
rect 10850 5414 10862 5466
rect 10924 5414 10926 5466
rect 10764 5412 10788 5414
rect 10844 5412 10868 5414
rect 10924 5412 10948 5414
rect 10708 5392 11004 5412
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10598 4992 10654 5001
rect 10598 4927 10654 4936
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10232 4548 10284 4554
rect 10232 4490 10284 4496
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10152 4146 10180 4422
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10152 3534 10180 4082
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 9404 2440 9456 2446
rect 9232 2378 9352 2394
rect 9404 2382 9456 2388
rect 9036 2372 9088 2378
rect 9232 2372 9364 2378
rect 9232 2366 9312 2372
rect 9036 2314 9088 2320
rect 9312 2314 9364 2320
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9232 800 9260 2246
rect 10244 2106 10272 2314
rect 10232 2100 10284 2106
rect 10232 2042 10284 2048
rect 10520 1154 10548 4626
rect 10612 1970 10640 4927
rect 11072 4826 11100 6326
rect 11164 6254 11192 7142
rect 11348 6390 11376 7686
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11072 4622 11100 4762
rect 11060 4616 11112 4622
rect 11440 4593 11468 8910
rect 11532 8498 11560 10406
rect 11624 9489 11652 13892
rect 11704 13874 11756 13880
rect 11900 13394 12020 13410
rect 11888 13388 12020 13394
rect 11940 13382 12020 13388
rect 11888 13330 11940 13336
rect 11888 13252 11940 13258
rect 11888 13194 11940 13200
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11716 12238 11744 12786
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11716 11626 11744 12174
rect 11808 12102 11836 12582
rect 11900 12442 11928 13194
rect 11992 12850 12020 13382
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11796 12096 11848 12102
rect 11980 12096 12032 12102
rect 11848 12044 11928 12050
rect 11796 12038 11928 12044
rect 11980 12038 12032 12044
rect 11808 12022 11928 12038
rect 11808 11973 11836 12022
rect 11900 11762 11928 12022
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11704 11620 11756 11626
rect 11704 11562 11756 11568
rect 11992 11558 12020 12038
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11992 11354 12020 11494
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11900 10266 11928 11086
rect 12084 10810 12112 14350
rect 12176 13394 12204 14350
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12176 13258 12204 13330
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12176 11150 12204 12786
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11716 9518 11744 9998
rect 11900 9994 11928 10066
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11808 9722 11836 9930
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11808 9586 11836 9658
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11704 9512 11756 9518
rect 11610 9480 11666 9489
rect 11900 9466 11928 9590
rect 11704 9454 11756 9460
rect 11610 9415 11666 9424
rect 11808 9438 11928 9466
rect 11808 9364 11836 9438
rect 11624 9336 11836 9364
rect 11624 8974 11652 9336
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11992 8922 12020 10678
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12084 10044 12112 10610
rect 12176 10266 12204 11086
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12164 10056 12216 10062
rect 12084 10024 12164 10044
rect 12216 10024 12218 10033
rect 12084 10016 12162 10024
rect 12162 9959 12218 9968
rect 12268 9382 12296 13874
rect 12452 13326 12480 14486
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12636 13818 12664 14418
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12728 14006 12756 14350
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12820 13938 12848 14350
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12912 13818 12940 14878
rect 12544 13530 12572 13806
rect 12636 13790 12756 13818
rect 12820 13802 12940 13818
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 12170 12480 12582
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12360 9518 12388 11154
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12452 10198 12480 11018
rect 12636 10690 12664 13670
rect 12728 11354 12756 13790
rect 12808 13796 12940 13802
rect 12860 13790 12940 13796
rect 12808 13738 12860 13744
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12912 12306 12940 13262
rect 13004 12628 13032 15438
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13146 14716 13442 14736
rect 13202 14714 13226 14716
rect 13282 14714 13306 14716
rect 13362 14714 13386 14716
rect 13224 14662 13226 14714
rect 13288 14662 13300 14714
rect 13362 14662 13364 14714
rect 13202 14660 13226 14662
rect 13282 14660 13306 14662
rect 13362 14660 13386 14662
rect 13146 14640 13442 14660
rect 13556 14618 13584 14894
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13740 14482 13768 14894
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13146 13628 13442 13648
rect 13202 13626 13226 13628
rect 13282 13626 13306 13628
rect 13362 13626 13386 13628
rect 13224 13574 13226 13626
rect 13288 13574 13300 13626
rect 13362 13574 13364 13626
rect 13202 13572 13226 13574
rect 13282 13572 13306 13574
rect 13362 13572 13386 13574
rect 13146 13552 13442 13572
rect 13556 13530 13584 13806
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13648 13326 13676 13738
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13740 12918 13768 14418
rect 13832 13938 13860 15914
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13924 14550 13952 14894
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 13924 14074 13952 14486
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13728 12912 13780 12918
rect 13728 12854 13780 12860
rect 13004 12600 13584 12628
rect 13146 12540 13442 12560
rect 13202 12538 13226 12540
rect 13282 12538 13306 12540
rect 13362 12538 13386 12540
rect 13224 12486 13226 12538
rect 13288 12486 13300 12538
rect 13362 12486 13364 12538
rect 13202 12484 13226 12486
rect 13282 12484 13306 12486
rect 13362 12484 13386 12486
rect 13146 12464 13442 12484
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12912 11830 12940 12038
rect 12900 11824 12952 11830
rect 12900 11766 12952 11772
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12820 11286 12848 11630
rect 12912 11354 12940 11766
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 13004 11150 13032 11494
rect 13146 11452 13442 11472
rect 13202 11450 13226 11452
rect 13282 11450 13306 11452
rect 13362 11450 13386 11452
rect 13224 11398 13226 11450
rect 13288 11398 13300 11450
rect 13362 11398 13364 11450
rect 13202 11396 13226 11398
rect 13282 11396 13306 11398
rect 13362 11396 13386 11398
rect 13146 11376 13442 11396
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12912 10962 12940 11086
rect 13096 10962 13124 11222
rect 12912 10934 13124 10962
rect 12544 10662 12664 10690
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 12716 10668 12768 10674
rect 12440 10192 12492 10198
rect 12438 10160 12440 10169
rect 12492 10160 12494 10169
rect 12438 10095 12494 10104
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12452 9722 12480 9998
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11624 8430 11652 8910
rect 11992 8894 12112 8922
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11624 7818 11652 8366
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11612 7812 11664 7818
rect 11612 7754 11664 7760
rect 11716 7750 11744 7890
rect 11900 7886 11928 8366
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11624 6254 11652 6938
rect 11716 6458 11744 7686
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11808 6458 11836 7346
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11808 6322 11836 6394
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11624 5370 11744 5386
rect 11612 5364 11744 5370
rect 11664 5358 11744 5364
rect 11612 5306 11664 5312
rect 11520 5296 11572 5302
rect 11518 5264 11520 5273
rect 11572 5264 11574 5273
rect 11518 5199 11574 5208
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11610 5128 11666 5137
rect 11532 4622 11560 5102
rect 11610 5063 11666 5072
rect 11520 4616 11572 4622
rect 11060 4558 11112 4564
rect 11426 4584 11482 4593
rect 11520 4558 11572 4564
rect 11624 4554 11652 5063
rect 11426 4519 11482 4528
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10708 4380 11004 4400
rect 10764 4378 10788 4380
rect 10844 4378 10868 4380
rect 10924 4378 10948 4380
rect 10786 4326 10788 4378
rect 10850 4326 10862 4378
rect 10924 4326 10926 4378
rect 10764 4324 10788 4326
rect 10844 4324 10868 4326
rect 10924 4324 10948 4326
rect 10708 4304 11004 4324
rect 11072 3534 11100 4422
rect 11716 4146 11744 5358
rect 11808 5234 11836 5510
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11808 4690 11836 5170
rect 11900 4758 11928 7414
rect 11992 7342 12020 8774
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11992 7002 12020 7278
rect 12084 7206 12112 8894
rect 12452 7993 12480 9046
rect 12438 7984 12494 7993
rect 12438 7919 12494 7928
rect 12544 7818 12572 10662
rect 12716 10610 12768 10616
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12544 7478 12572 7754
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12452 7206 12480 7346
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 12084 6644 12112 7142
rect 12268 6798 12296 7142
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12164 6656 12216 6662
rect 12084 6616 12164 6644
rect 12164 6598 12216 6604
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11992 5846 12020 6258
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 12070 5808 12126 5817
rect 12070 5743 12126 5752
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11992 5137 12020 5170
rect 11978 5128 12034 5137
rect 11978 5063 12034 5072
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11900 4078 11928 4558
rect 12084 4434 12112 5743
rect 12176 5234 12204 6054
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 11992 4406 12112 4434
rect 11992 4146 12020 4406
rect 12268 4264 12296 6054
rect 12360 5710 12388 6938
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12438 5264 12494 5273
rect 12438 5199 12440 5208
rect 12492 5199 12494 5208
rect 12440 5170 12492 5176
rect 12452 5030 12480 5170
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12544 4758 12572 7210
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12084 4236 12296 4264
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11256 3534 11284 3878
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 10708 3292 11004 3312
rect 10764 3290 10788 3292
rect 10844 3290 10868 3292
rect 10924 3290 10948 3292
rect 10786 3238 10788 3290
rect 10850 3238 10862 3290
rect 10924 3238 10926 3290
rect 10764 3236 10788 3238
rect 10844 3236 10868 3238
rect 10924 3236 10948 3238
rect 10708 3216 11004 3236
rect 11072 3058 11100 3470
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 3194 11192 3402
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 11164 2650 11192 2858
rect 11256 2650 11284 3470
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11532 2446 11560 3130
rect 11808 3126 11836 3334
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11808 2446 11836 3062
rect 11900 3058 11928 3470
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 11992 2990 12020 3946
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 11992 2446 12020 2926
rect 12084 2854 12112 4236
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 12162 2952 12218 2961
rect 12268 2922 12296 3470
rect 12162 2887 12218 2896
rect 12256 2916 12308 2922
rect 12176 2854 12204 2887
rect 12256 2858 12308 2864
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 12544 2650 12572 4422
rect 12636 4146 12664 10542
rect 12728 8294 12756 10610
rect 13096 10538 13124 10678
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13146 10364 13442 10384
rect 13202 10362 13226 10364
rect 13282 10362 13306 10364
rect 13362 10362 13386 10364
rect 13224 10310 13226 10362
rect 13288 10310 13300 10362
rect 13362 10310 13364 10362
rect 13202 10308 13226 10310
rect 13282 10308 13306 10310
rect 13362 10308 13386 10310
rect 13146 10288 13442 10308
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13004 10010 13032 10202
rect 13084 10192 13136 10198
rect 13082 10160 13084 10169
rect 13136 10160 13138 10169
rect 13082 10095 13138 10104
rect 13268 10056 13320 10062
rect 13004 9982 13124 10010
rect 13268 9998 13320 10004
rect 13358 10024 13414 10033
rect 13096 9926 13124 9982
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13280 9722 13308 9998
rect 13358 9959 13360 9968
rect 13412 9959 13414 9968
rect 13360 9930 13412 9936
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 12820 9586 12848 9658
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 9178 12848 9522
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12912 8498 12940 9454
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 13004 8566 13032 9318
rect 13146 9276 13442 9296
rect 13202 9274 13226 9276
rect 13282 9274 13306 9276
rect 13362 9274 13386 9276
rect 13224 9222 13226 9274
rect 13288 9222 13300 9274
rect 13362 9222 13364 9274
rect 13202 9220 13226 9222
rect 13282 9220 13306 9222
rect 13362 9220 13386 9222
rect 13146 9200 13442 9220
rect 13556 9058 13584 12600
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 13464 9030 13584 9058
rect 12992 8560 13044 8566
rect 12992 8502 13044 8508
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12728 7886 12756 8230
rect 12820 8129 12848 8366
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12806 8120 12862 8129
rect 12806 8055 12862 8064
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12912 7478 12940 8230
rect 13004 7970 13032 8502
rect 13464 8430 13492 9030
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13146 8188 13442 8208
rect 13202 8186 13226 8188
rect 13282 8186 13306 8188
rect 13362 8186 13386 8188
rect 13224 8134 13226 8186
rect 13288 8134 13300 8186
rect 13362 8134 13364 8186
rect 13202 8132 13226 8134
rect 13282 8132 13306 8134
rect 13362 8132 13386 8134
rect 13146 8112 13442 8132
rect 13004 7942 13124 7970
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12820 7002 12848 7142
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12912 6798 12940 7414
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 13004 6730 13032 7686
rect 13096 7410 13124 7942
rect 13556 7886 13584 8434
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13556 7546 13584 7822
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13146 7100 13442 7120
rect 13202 7098 13226 7100
rect 13282 7098 13306 7100
rect 13362 7098 13386 7100
rect 13224 7046 13226 7098
rect 13288 7046 13300 7098
rect 13362 7046 13364 7098
rect 13202 7044 13226 7046
rect 13282 7044 13306 7046
rect 13362 7044 13386 7046
rect 13146 7024 13442 7044
rect 13648 6914 13676 11222
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13740 10470 13768 10610
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10062 13768 10406
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13740 8634 13768 9522
rect 13832 9450 13860 11562
rect 13924 11354 13952 13806
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13924 10606 13952 10950
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13832 8974 13860 9386
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13740 7818 13768 8570
rect 13832 8022 13860 8910
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13556 6886 13676 6914
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 13004 6322 13032 6666
rect 12808 6316 12860 6322
rect 12992 6316 13044 6322
rect 12808 6258 12860 6264
rect 12912 6276 12992 6304
rect 12820 5914 12848 6258
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12806 5808 12862 5817
rect 12806 5743 12862 5752
rect 12820 5710 12848 5743
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12728 4282 12756 4626
rect 12820 4554 12848 5510
rect 12912 4729 12940 6276
rect 12992 6258 13044 6264
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 13004 5370 13032 6122
rect 13146 6012 13442 6032
rect 13202 6010 13226 6012
rect 13282 6010 13306 6012
rect 13362 6010 13386 6012
rect 13224 5958 13226 6010
rect 13288 5958 13300 6010
rect 13362 5958 13364 6010
rect 13202 5956 13226 5958
rect 13282 5956 13306 5958
rect 13362 5956 13386 5958
rect 13146 5936 13442 5956
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 13464 5234 13492 5646
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13004 4826 13032 5170
rect 13146 4924 13442 4944
rect 13202 4922 13226 4924
rect 13282 4922 13306 4924
rect 13362 4922 13386 4924
rect 13224 4870 13226 4922
rect 13288 4870 13300 4922
rect 13362 4870 13364 4922
rect 13202 4868 13226 4870
rect 13282 4868 13306 4870
rect 13362 4868 13386 4870
rect 13146 4848 13442 4868
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 12898 4720 12954 4729
rect 12898 4655 12954 4664
rect 12808 4548 12860 4554
rect 12808 4490 12860 4496
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12820 4214 12848 4490
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12624 4140 12676 4146
rect 12676 4100 12756 4128
rect 12624 4082 12676 4088
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12636 2446 12664 3674
rect 12728 3670 12756 4100
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12912 3602 12940 4218
rect 13004 4214 13032 4762
rect 13266 4720 13322 4729
rect 13556 4706 13584 6886
rect 13740 6866 13768 7754
rect 13832 7342 13860 7958
rect 13924 7342 13952 10542
rect 14016 8430 14044 15302
rect 14200 13546 14228 15438
rect 14292 14414 14320 15438
rect 14464 15428 14516 15434
rect 14464 15370 14516 15376
rect 14476 15162 14504 15370
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14476 14414 14504 15098
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14200 13518 14320 13546
rect 14188 13456 14240 13462
rect 14188 13398 14240 13404
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14108 12782 14136 13262
rect 14200 12782 14228 13398
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14200 12442 14228 12718
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 5166 13676 6734
rect 13832 6322 13860 7142
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13832 5710 13860 6258
rect 14016 5846 14044 8366
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13910 5672 13966 5681
rect 13910 5607 13966 5616
rect 13924 5302 13952 5607
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 13912 5296 13964 5302
rect 13912 5238 13964 5244
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13266 4655 13322 4664
rect 13464 4678 13584 4706
rect 13280 4622 13308 4655
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13096 4486 13124 4558
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 12992 4208 13044 4214
rect 12992 4150 13044 4156
rect 13372 4146 13400 4558
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13464 4010 13492 4678
rect 13544 4636 13596 4642
rect 13544 4578 13596 4584
rect 13728 4616 13780 4622
rect 13556 4078 13584 4578
rect 13728 4558 13780 4564
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13146 3836 13442 3856
rect 13202 3834 13226 3836
rect 13282 3834 13306 3836
rect 13362 3834 13386 3836
rect 13224 3782 13226 3834
rect 13288 3782 13300 3834
rect 13362 3782 13364 3834
rect 13202 3780 13226 3782
rect 13282 3780 13306 3782
rect 13362 3780 13386 3782
rect 13146 3760 13442 3780
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 12912 3058 12940 3538
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 13146 2748 13442 2768
rect 13202 2746 13226 2748
rect 13282 2746 13306 2748
rect 13362 2746 13386 2748
rect 13224 2694 13226 2746
rect 13288 2694 13300 2746
rect 13362 2694 13364 2746
rect 13202 2692 13226 2694
rect 13282 2692 13306 2694
rect 13362 2692 13386 2694
rect 13146 2672 13442 2692
rect 13556 2553 13584 3402
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 3058 13676 3334
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 13740 2582 13768 4558
rect 13912 4548 13964 4554
rect 13912 4490 13964 4496
rect 13924 4010 13952 4490
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13728 2576 13780 2582
rect 13542 2544 13598 2553
rect 13728 2518 13780 2524
rect 13542 2479 13598 2488
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 13924 2378 13952 3946
rect 14016 3534 14044 5510
rect 14108 3738 14136 11698
rect 14292 9518 14320 13518
rect 14384 10198 14412 14214
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14476 12986 14504 13262
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14476 12102 14504 12922
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14568 11218 14596 16050
rect 14660 15706 14688 16050
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14752 14498 14780 15846
rect 14936 15366 14964 18215
rect 16776 16182 16804 18215
rect 16764 16176 16816 16182
rect 15014 16144 15070 16153
rect 16764 16118 16816 16124
rect 15014 16079 15016 16088
rect 15068 16079 15070 16088
rect 15016 16050 15068 16056
rect 14924 15360 14976 15366
rect 14924 15302 14976 15308
rect 14660 14470 14780 14498
rect 14660 13410 14688 14470
rect 14740 14340 14792 14346
rect 14740 14282 14792 14288
rect 14752 13530 14780 14282
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14660 13382 14780 13410
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14660 12374 14688 13262
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14752 11354 14780 13382
rect 14844 12442 14872 13874
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15028 13433 15056 13806
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 15014 13424 15070 13433
rect 15014 13359 15070 13368
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14292 8498 14320 9454
rect 14384 8974 14412 10134
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14476 9178 14504 9454
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14476 8634 14504 9114
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14568 8362 14596 11154
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14200 5370 14228 7346
rect 14292 6458 14320 7822
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14384 6866 14412 7278
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14292 6338 14320 6394
rect 14292 6310 14412 6338
rect 14280 5840 14332 5846
rect 14280 5782 14332 5788
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14292 5234 14320 5782
rect 14384 5778 14412 6310
rect 14476 5914 14504 7346
rect 14660 6746 14688 10610
rect 14740 10532 14792 10538
rect 14740 10474 14792 10480
rect 14568 6718 14688 6746
rect 14568 6254 14596 6718
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14568 5778 14596 6190
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4758 14228 4966
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14200 4146 14228 4694
rect 14476 4690 14504 5034
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14568 4622 14596 5578
rect 14660 4758 14688 6598
rect 14648 4752 14700 4758
rect 14648 4694 14700 4700
rect 14556 4616 14608 4622
rect 14462 4584 14518 4593
rect 14556 4558 14608 4564
rect 14462 4519 14518 4528
rect 14476 4282 14504 4519
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14292 3534 14320 4082
rect 14476 3602 14504 4218
rect 14660 4146 14688 4694
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14660 2990 14688 3470
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14660 2650 14688 2926
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 14372 2576 14424 2582
rect 14372 2518 14424 2524
rect 14384 2378 14412 2518
rect 14752 2446 14780 10474
rect 14844 9602 14872 11630
rect 14936 10713 14964 11698
rect 14922 10704 14978 10713
rect 14922 10639 14978 10648
rect 14844 9574 14964 9602
rect 15120 9586 15148 13670
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14844 8362 14872 9454
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14844 5642 14872 6054
rect 14936 5642 14964 9574
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15120 9194 15148 9522
rect 15120 9166 15240 9194
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 14832 5636 14884 5642
rect 14832 5578 14884 5584
rect 14924 5636 14976 5642
rect 14924 5578 14976 5584
rect 15028 5522 15056 8842
rect 15212 8634 15240 9166
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 14844 5494 15056 5522
rect 14844 2582 14872 5494
rect 15014 5264 15070 5273
rect 15014 5199 15016 5208
rect 15068 5199 15070 5208
rect 15016 5170 15068 5176
rect 14832 2576 14884 2582
rect 14832 2518 14884 2524
rect 14844 2446 14872 2518
rect 14924 2508 14976 2514
rect 14924 2450 14976 2456
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 13912 2372 13964 2378
rect 13912 2314 13964 2320
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 14752 2310 14780 2382
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 10708 2204 11004 2224
rect 10764 2202 10788 2204
rect 10844 2202 10868 2204
rect 10924 2202 10948 2204
rect 10786 2150 10788 2202
rect 10850 2150 10862 2202
rect 10924 2150 10926 2202
rect 10764 2148 10788 2150
rect 10844 2148 10868 2150
rect 10924 2148 10948 2150
rect 10708 2128 11004 2148
rect 10600 1964 10652 1970
rect 10600 1906 10652 1912
rect 12900 1964 12952 1970
rect 12900 1906 12952 1912
rect 10508 1148 10560 1154
rect 10508 1090 10560 1096
rect 11060 1148 11112 1154
rect 11060 1090 11112 1096
rect 11072 800 11100 1090
rect 12912 800 12940 1906
rect 14936 800 14964 2450
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 16776 800 16804 2314
rect 18 0 74 800
rect 1858 0 1914 800
rect 3698 0 3754 800
rect 5538 0 5594 800
rect 7378 0 7434 800
rect 9218 0 9274 800
rect 11058 0 11114 800
rect 12898 0 12954 800
rect 14922 0 14978 800
rect 16762 0 16818 800
<< via2 >>
rect 1398 16360 1454 16416
rect 5832 16346 5888 16348
rect 5912 16346 5968 16348
rect 5992 16346 6048 16348
rect 6072 16346 6128 16348
rect 5832 16294 5858 16346
rect 5858 16294 5888 16346
rect 5912 16294 5922 16346
rect 5922 16294 5968 16346
rect 5992 16294 6038 16346
rect 6038 16294 6048 16346
rect 6072 16294 6102 16346
rect 6102 16294 6128 16346
rect 5832 16292 5888 16294
rect 5912 16292 5968 16294
rect 5992 16292 6048 16294
rect 6072 16292 6128 16294
rect 10708 16346 10764 16348
rect 10788 16346 10844 16348
rect 10868 16346 10924 16348
rect 10948 16346 11004 16348
rect 10708 16294 10734 16346
rect 10734 16294 10764 16346
rect 10788 16294 10798 16346
rect 10798 16294 10844 16346
rect 10868 16294 10914 16346
rect 10914 16294 10924 16346
rect 10948 16294 10978 16346
rect 10978 16294 11004 16346
rect 10708 16292 10764 16294
rect 10788 16292 10844 16294
rect 10868 16292 10924 16294
rect 10948 16292 11004 16294
rect 1858 13640 1914 13696
rect 1858 10920 1914 10976
rect 3394 15802 3450 15804
rect 3474 15802 3530 15804
rect 3554 15802 3610 15804
rect 3634 15802 3690 15804
rect 3394 15750 3420 15802
rect 3420 15750 3450 15802
rect 3474 15750 3484 15802
rect 3484 15750 3530 15802
rect 3554 15750 3600 15802
rect 3600 15750 3610 15802
rect 3634 15750 3664 15802
rect 3664 15750 3690 15802
rect 3394 15748 3450 15750
rect 3474 15748 3530 15750
rect 3554 15748 3610 15750
rect 3634 15748 3690 15750
rect 3394 14714 3450 14716
rect 3474 14714 3530 14716
rect 3554 14714 3610 14716
rect 3634 14714 3690 14716
rect 3394 14662 3420 14714
rect 3420 14662 3450 14714
rect 3474 14662 3484 14714
rect 3484 14662 3530 14714
rect 3554 14662 3600 14714
rect 3600 14662 3610 14714
rect 3634 14662 3664 14714
rect 3664 14662 3690 14714
rect 3394 14660 3450 14662
rect 3474 14660 3530 14662
rect 3554 14660 3610 14662
rect 3634 14660 3690 14662
rect 3394 13626 3450 13628
rect 3474 13626 3530 13628
rect 3554 13626 3610 13628
rect 3634 13626 3690 13628
rect 3394 13574 3420 13626
rect 3420 13574 3450 13626
rect 3474 13574 3484 13626
rect 3484 13574 3530 13626
rect 3554 13574 3600 13626
rect 3600 13574 3610 13626
rect 3634 13574 3664 13626
rect 3664 13574 3690 13626
rect 3394 13572 3450 13574
rect 3474 13572 3530 13574
rect 3554 13572 3610 13574
rect 3634 13572 3690 13574
rect 3394 12538 3450 12540
rect 3474 12538 3530 12540
rect 3554 12538 3610 12540
rect 3634 12538 3690 12540
rect 3394 12486 3420 12538
rect 3420 12486 3450 12538
rect 3474 12486 3484 12538
rect 3484 12486 3530 12538
rect 3554 12486 3600 12538
rect 3600 12486 3610 12538
rect 3634 12486 3664 12538
rect 3664 12486 3690 12538
rect 3394 12484 3450 12486
rect 3474 12484 3530 12486
rect 3554 12484 3610 12486
rect 3634 12484 3690 12486
rect 3394 11450 3450 11452
rect 3474 11450 3530 11452
rect 3554 11450 3610 11452
rect 3634 11450 3690 11452
rect 3394 11398 3420 11450
rect 3420 11398 3450 11450
rect 3474 11398 3484 11450
rect 3484 11398 3530 11450
rect 3554 11398 3600 11450
rect 3600 11398 3610 11450
rect 3634 11398 3664 11450
rect 3664 11398 3690 11450
rect 3394 11396 3450 11398
rect 3474 11396 3530 11398
rect 3554 11396 3610 11398
rect 3634 11396 3690 11398
rect 3394 10362 3450 10364
rect 3474 10362 3530 10364
rect 3554 10362 3610 10364
rect 3634 10362 3690 10364
rect 3394 10310 3420 10362
rect 3420 10310 3450 10362
rect 3474 10310 3484 10362
rect 3484 10310 3530 10362
rect 3554 10310 3600 10362
rect 3600 10310 3610 10362
rect 3634 10310 3664 10362
rect 3664 10310 3690 10362
rect 3394 10308 3450 10310
rect 3474 10308 3530 10310
rect 3554 10308 3610 10310
rect 3634 10308 3690 10310
rect 3790 9424 3846 9480
rect 3394 9274 3450 9276
rect 3474 9274 3530 9276
rect 3554 9274 3610 9276
rect 3634 9274 3690 9276
rect 3394 9222 3420 9274
rect 3420 9222 3450 9274
rect 3474 9222 3484 9274
rect 3484 9222 3530 9274
rect 3554 9222 3600 9274
rect 3600 9222 3610 9274
rect 3634 9222 3664 9274
rect 3664 9222 3690 9274
rect 3394 9220 3450 9222
rect 3474 9220 3530 9222
rect 3554 9220 3610 9222
rect 3634 9220 3690 9222
rect 2870 8200 2926 8256
rect 3394 8186 3450 8188
rect 3474 8186 3530 8188
rect 3554 8186 3610 8188
rect 3634 8186 3690 8188
rect 3394 8134 3420 8186
rect 3420 8134 3450 8186
rect 3474 8134 3484 8186
rect 3484 8134 3530 8186
rect 3554 8134 3600 8186
rect 3600 8134 3610 8186
rect 3634 8134 3664 8186
rect 3664 8134 3690 8186
rect 3394 8132 3450 8134
rect 3474 8132 3530 8134
rect 3554 8132 3610 8134
rect 3634 8132 3690 8134
rect 2410 5652 2412 5672
rect 2412 5652 2464 5672
rect 2464 5652 2466 5672
rect 2410 5616 2466 5652
rect 1398 5480 1454 5536
rect 3394 7098 3450 7100
rect 3474 7098 3530 7100
rect 3554 7098 3610 7100
rect 3634 7098 3690 7100
rect 3394 7046 3420 7098
rect 3420 7046 3450 7098
rect 3474 7046 3484 7098
rect 3484 7046 3530 7098
rect 3554 7046 3600 7098
rect 3600 7046 3610 7098
rect 3634 7046 3664 7098
rect 3664 7046 3690 7098
rect 3394 7044 3450 7046
rect 3474 7044 3530 7046
rect 3554 7044 3610 7046
rect 3634 7044 3690 7046
rect 2410 5072 2466 5128
rect 3394 6010 3450 6012
rect 3474 6010 3530 6012
rect 3554 6010 3610 6012
rect 3634 6010 3690 6012
rect 3394 5958 3420 6010
rect 3420 5958 3450 6010
rect 3474 5958 3484 6010
rect 3484 5958 3530 6010
rect 3554 5958 3600 6010
rect 3600 5958 3610 6010
rect 3634 5958 3664 6010
rect 3664 5958 3690 6010
rect 3394 5956 3450 5958
rect 3474 5956 3530 5958
rect 3554 5956 3610 5958
rect 3634 5956 3690 5958
rect 5832 15258 5888 15260
rect 5912 15258 5968 15260
rect 5992 15258 6048 15260
rect 6072 15258 6128 15260
rect 5832 15206 5858 15258
rect 5858 15206 5888 15258
rect 5912 15206 5922 15258
rect 5922 15206 5968 15258
rect 5992 15206 6038 15258
rect 6038 15206 6048 15258
rect 6072 15206 6102 15258
rect 6102 15206 6128 15258
rect 5832 15204 5888 15206
rect 5912 15204 5968 15206
rect 5992 15204 6048 15206
rect 6072 15204 6128 15206
rect 5832 14170 5888 14172
rect 5912 14170 5968 14172
rect 5992 14170 6048 14172
rect 6072 14170 6128 14172
rect 5832 14118 5858 14170
rect 5858 14118 5888 14170
rect 5912 14118 5922 14170
rect 5922 14118 5968 14170
rect 5992 14118 6038 14170
rect 6038 14118 6048 14170
rect 6072 14118 6102 14170
rect 6102 14118 6128 14170
rect 5832 14116 5888 14118
rect 5912 14116 5968 14118
rect 5992 14116 6048 14118
rect 6072 14116 6128 14118
rect 5832 13082 5888 13084
rect 5912 13082 5968 13084
rect 5992 13082 6048 13084
rect 6072 13082 6128 13084
rect 5832 13030 5858 13082
rect 5858 13030 5888 13082
rect 5912 13030 5922 13082
rect 5922 13030 5968 13082
rect 5992 13030 6038 13082
rect 6038 13030 6048 13082
rect 6072 13030 6102 13082
rect 6102 13030 6128 13082
rect 5832 13028 5888 13030
rect 5912 13028 5968 13030
rect 5992 13028 6048 13030
rect 6072 13028 6128 13030
rect 3394 4922 3450 4924
rect 3474 4922 3530 4924
rect 3554 4922 3610 4924
rect 3634 4922 3690 4924
rect 3394 4870 3420 4922
rect 3420 4870 3450 4922
rect 3474 4870 3484 4922
rect 3484 4870 3530 4922
rect 3554 4870 3600 4922
rect 3600 4870 3610 4922
rect 3634 4870 3664 4922
rect 3664 4870 3690 4922
rect 3394 4868 3450 4870
rect 3474 4868 3530 4870
rect 3554 4868 3610 4870
rect 3634 4868 3690 4870
rect 1398 2760 1454 2816
rect 3394 3834 3450 3836
rect 3474 3834 3530 3836
rect 3554 3834 3610 3836
rect 3634 3834 3690 3836
rect 3394 3782 3420 3834
rect 3420 3782 3450 3834
rect 3474 3782 3484 3834
rect 3484 3782 3530 3834
rect 3554 3782 3600 3834
rect 3600 3782 3610 3834
rect 3634 3782 3664 3834
rect 3664 3782 3690 3834
rect 3394 3780 3450 3782
rect 3474 3780 3530 3782
rect 3554 3780 3610 3782
rect 3634 3780 3690 3782
rect 5832 11994 5888 11996
rect 5912 11994 5968 11996
rect 5992 11994 6048 11996
rect 6072 11994 6128 11996
rect 5832 11942 5858 11994
rect 5858 11942 5888 11994
rect 5912 11942 5922 11994
rect 5922 11942 5968 11994
rect 5992 11942 6038 11994
rect 6038 11942 6048 11994
rect 6072 11942 6102 11994
rect 6102 11942 6128 11994
rect 5832 11940 5888 11942
rect 5912 11940 5968 11942
rect 5992 11940 6048 11942
rect 6072 11940 6128 11942
rect 5832 10906 5888 10908
rect 5912 10906 5968 10908
rect 5992 10906 6048 10908
rect 6072 10906 6128 10908
rect 5832 10854 5858 10906
rect 5858 10854 5888 10906
rect 5912 10854 5922 10906
rect 5922 10854 5968 10906
rect 5992 10854 6038 10906
rect 6038 10854 6048 10906
rect 6072 10854 6102 10906
rect 6102 10854 6128 10906
rect 5832 10852 5888 10854
rect 5912 10852 5968 10854
rect 5992 10852 6048 10854
rect 6072 10852 6128 10854
rect 5722 10668 5778 10704
rect 5722 10648 5724 10668
rect 5724 10648 5776 10668
rect 5776 10648 5778 10668
rect 5832 9818 5888 9820
rect 5912 9818 5968 9820
rect 5992 9818 6048 9820
rect 6072 9818 6128 9820
rect 5832 9766 5858 9818
rect 5858 9766 5888 9818
rect 5912 9766 5922 9818
rect 5922 9766 5968 9818
rect 5992 9766 6038 9818
rect 6038 9766 6048 9818
rect 6072 9766 6102 9818
rect 6102 9766 6128 9818
rect 5832 9764 5888 9766
rect 5912 9764 5968 9766
rect 5992 9764 6048 9766
rect 6072 9764 6128 9766
rect 5630 9580 5686 9616
rect 5630 9560 5632 9580
rect 5632 9560 5684 9580
rect 5684 9560 5686 9580
rect 5722 9424 5778 9480
rect 5832 8730 5888 8732
rect 5912 8730 5968 8732
rect 5992 8730 6048 8732
rect 6072 8730 6128 8732
rect 5832 8678 5858 8730
rect 5858 8678 5888 8730
rect 5912 8678 5922 8730
rect 5922 8678 5968 8730
rect 5992 8678 6038 8730
rect 6038 8678 6048 8730
rect 6072 8678 6102 8730
rect 6102 8678 6128 8730
rect 5832 8676 5888 8678
rect 5912 8676 5968 8678
rect 5992 8676 6048 8678
rect 6072 8676 6128 8678
rect 5832 7642 5888 7644
rect 5912 7642 5968 7644
rect 5992 7642 6048 7644
rect 6072 7642 6128 7644
rect 5832 7590 5858 7642
rect 5858 7590 5888 7642
rect 5912 7590 5922 7642
rect 5922 7590 5968 7642
rect 5992 7590 6038 7642
rect 6038 7590 6048 7642
rect 6072 7590 6102 7642
rect 6102 7590 6128 7642
rect 5832 7588 5888 7590
rect 5912 7588 5968 7590
rect 5992 7588 6048 7590
rect 6072 7588 6128 7590
rect 5832 6554 5888 6556
rect 5912 6554 5968 6556
rect 5992 6554 6048 6556
rect 6072 6554 6128 6556
rect 5832 6502 5858 6554
rect 5858 6502 5888 6554
rect 5912 6502 5922 6554
rect 5922 6502 5968 6554
rect 5992 6502 6038 6554
rect 6038 6502 6048 6554
rect 6072 6502 6102 6554
rect 6102 6502 6128 6554
rect 5832 6500 5888 6502
rect 5912 6500 5968 6502
rect 5992 6500 6048 6502
rect 6072 6500 6128 6502
rect 3394 2746 3450 2748
rect 3474 2746 3530 2748
rect 3554 2746 3610 2748
rect 3634 2746 3690 2748
rect 3394 2694 3420 2746
rect 3420 2694 3450 2746
rect 3474 2694 3484 2746
rect 3484 2694 3530 2746
rect 3554 2694 3600 2746
rect 3600 2694 3610 2746
rect 3634 2694 3664 2746
rect 3664 2694 3690 2746
rect 3394 2692 3450 2694
rect 3474 2692 3530 2694
rect 3554 2692 3610 2694
rect 3634 2692 3690 2694
rect 5832 5466 5888 5468
rect 5912 5466 5968 5468
rect 5992 5466 6048 5468
rect 6072 5466 6128 5468
rect 5832 5414 5858 5466
rect 5858 5414 5888 5466
rect 5912 5414 5922 5466
rect 5922 5414 5968 5466
rect 5992 5414 6038 5466
rect 6038 5414 6048 5466
rect 6072 5414 6102 5466
rect 6102 5414 6128 5466
rect 5832 5412 5888 5414
rect 5912 5412 5968 5414
rect 5992 5412 6048 5414
rect 6072 5412 6128 5414
rect 6182 5208 6238 5264
rect 5832 4378 5888 4380
rect 5912 4378 5968 4380
rect 5992 4378 6048 4380
rect 6072 4378 6128 4380
rect 5832 4326 5858 4378
rect 5858 4326 5888 4378
rect 5912 4326 5922 4378
rect 5922 4326 5968 4378
rect 5992 4326 6038 4378
rect 6038 4326 6048 4378
rect 6072 4326 6102 4378
rect 6102 4326 6128 4378
rect 5832 4324 5888 4326
rect 5912 4324 5968 4326
rect 5992 4324 6048 4326
rect 6072 4324 6128 4326
rect 6274 4392 6330 4448
rect 5832 3290 5888 3292
rect 5912 3290 5968 3292
rect 5992 3290 6048 3292
rect 6072 3290 6128 3292
rect 5832 3238 5858 3290
rect 5858 3238 5888 3290
rect 5912 3238 5922 3290
rect 5922 3238 5968 3290
rect 5992 3238 6038 3290
rect 6038 3238 6048 3290
rect 6072 3238 6102 3290
rect 6102 3238 6128 3290
rect 5832 3236 5888 3238
rect 5912 3236 5968 3238
rect 5992 3236 6048 3238
rect 6072 3236 6128 3238
rect 5832 2202 5888 2204
rect 5912 2202 5968 2204
rect 5992 2202 6048 2204
rect 6072 2202 6128 2204
rect 5832 2150 5858 2202
rect 5858 2150 5888 2202
rect 5912 2150 5922 2202
rect 5922 2150 5968 2202
rect 5992 2150 6038 2202
rect 6038 2150 6048 2202
rect 6072 2150 6102 2202
rect 6102 2150 6128 2202
rect 5832 2148 5888 2150
rect 5912 2148 5968 2150
rect 5992 2148 6048 2150
rect 6072 2148 6128 2150
rect 8270 15802 8326 15804
rect 8350 15802 8406 15804
rect 8430 15802 8486 15804
rect 8510 15802 8566 15804
rect 8270 15750 8296 15802
rect 8296 15750 8326 15802
rect 8350 15750 8360 15802
rect 8360 15750 8406 15802
rect 8430 15750 8476 15802
rect 8476 15750 8486 15802
rect 8510 15750 8540 15802
rect 8540 15750 8566 15802
rect 8270 15748 8326 15750
rect 8350 15748 8406 15750
rect 8430 15748 8486 15750
rect 8510 15748 8566 15750
rect 8270 14714 8326 14716
rect 8350 14714 8406 14716
rect 8430 14714 8486 14716
rect 8510 14714 8566 14716
rect 8270 14662 8296 14714
rect 8296 14662 8326 14714
rect 8350 14662 8360 14714
rect 8360 14662 8406 14714
rect 8430 14662 8476 14714
rect 8476 14662 8486 14714
rect 8510 14662 8540 14714
rect 8540 14662 8566 14714
rect 8270 14660 8326 14662
rect 8350 14660 8406 14662
rect 8430 14660 8486 14662
rect 8510 14660 8566 14662
rect 7194 10668 7250 10704
rect 7194 10648 7196 10668
rect 7196 10648 7248 10668
rect 7248 10648 7250 10668
rect 7102 6432 7158 6488
rect 8270 13626 8326 13628
rect 8350 13626 8406 13628
rect 8430 13626 8486 13628
rect 8510 13626 8566 13628
rect 8270 13574 8296 13626
rect 8296 13574 8326 13626
rect 8350 13574 8360 13626
rect 8360 13574 8406 13626
rect 8430 13574 8476 13626
rect 8476 13574 8486 13626
rect 8510 13574 8540 13626
rect 8540 13574 8566 13626
rect 8270 13572 8326 13574
rect 8350 13572 8406 13574
rect 8430 13572 8486 13574
rect 8510 13572 8566 13574
rect 8270 12538 8326 12540
rect 8350 12538 8406 12540
rect 8430 12538 8486 12540
rect 8510 12538 8566 12540
rect 8270 12486 8296 12538
rect 8296 12486 8326 12538
rect 8350 12486 8360 12538
rect 8360 12486 8406 12538
rect 8430 12486 8476 12538
rect 8476 12486 8486 12538
rect 8510 12486 8540 12538
rect 8540 12486 8566 12538
rect 8270 12484 8326 12486
rect 8350 12484 8406 12486
rect 8430 12484 8486 12486
rect 8510 12484 8566 12486
rect 8270 11450 8326 11452
rect 8350 11450 8406 11452
rect 8430 11450 8486 11452
rect 8510 11450 8566 11452
rect 8270 11398 8296 11450
rect 8296 11398 8326 11450
rect 8350 11398 8360 11450
rect 8360 11398 8406 11450
rect 8430 11398 8476 11450
rect 8476 11398 8486 11450
rect 8510 11398 8540 11450
rect 8540 11398 8566 11450
rect 8270 11396 8326 11398
rect 8350 11396 8406 11398
rect 8430 11396 8486 11398
rect 8510 11396 8566 11398
rect 8270 10362 8326 10364
rect 8350 10362 8406 10364
rect 8430 10362 8486 10364
rect 8510 10362 8566 10364
rect 8270 10310 8296 10362
rect 8296 10310 8326 10362
rect 8350 10310 8360 10362
rect 8360 10310 8406 10362
rect 8430 10310 8476 10362
rect 8476 10310 8486 10362
rect 8510 10310 8540 10362
rect 8540 10310 8566 10362
rect 8270 10308 8326 10310
rect 8350 10308 8406 10310
rect 8430 10308 8486 10310
rect 8510 10308 8566 10310
rect 8114 9424 8170 9480
rect 8270 9274 8326 9276
rect 8350 9274 8406 9276
rect 8430 9274 8486 9276
rect 8510 9274 8566 9276
rect 8270 9222 8296 9274
rect 8296 9222 8326 9274
rect 8350 9222 8360 9274
rect 8360 9222 8406 9274
rect 8430 9222 8476 9274
rect 8476 9222 8486 9274
rect 8510 9222 8540 9274
rect 8540 9222 8566 9274
rect 8270 9220 8326 9222
rect 8350 9220 8406 9222
rect 8430 9220 8486 9222
rect 8510 9220 8566 9222
rect 8270 8186 8326 8188
rect 8350 8186 8406 8188
rect 8430 8186 8486 8188
rect 8510 8186 8566 8188
rect 8270 8134 8296 8186
rect 8296 8134 8326 8186
rect 8350 8134 8360 8186
rect 8360 8134 8406 8186
rect 8430 8134 8476 8186
rect 8476 8134 8486 8186
rect 8510 8134 8540 8186
rect 8540 8134 8566 8186
rect 8270 8132 8326 8134
rect 8350 8132 8406 8134
rect 8430 8132 8486 8134
rect 8510 8132 8566 8134
rect 8270 7098 8326 7100
rect 8350 7098 8406 7100
rect 8430 7098 8486 7100
rect 8510 7098 8566 7100
rect 8270 7046 8296 7098
rect 8296 7046 8326 7098
rect 8350 7046 8360 7098
rect 8360 7046 8406 7098
rect 8430 7046 8476 7098
rect 8476 7046 8486 7098
rect 8510 7046 8540 7098
rect 8540 7046 8566 7098
rect 8270 7044 8326 7046
rect 8350 7044 8406 7046
rect 8430 7044 8486 7046
rect 8510 7044 8566 7046
rect 7194 6316 7250 6352
rect 7194 6296 7196 6316
rect 7196 6296 7248 6316
rect 7248 6296 7250 6316
rect 6826 4528 6882 4584
rect 8574 6568 8630 6624
rect 8390 6160 8446 6216
rect 8270 6010 8326 6012
rect 8350 6010 8406 6012
rect 8430 6010 8486 6012
rect 8510 6010 8566 6012
rect 8270 5958 8296 6010
rect 8296 5958 8326 6010
rect 8350 5958 8360 6010
rect 8360 5958 8406 6010
rect 8430 5958 8476 6010
rect 8476 5958 8486 6010
rect 8510 5958 8540 6010
rect 8540 5958 8566 6010
rect 8270 5956 8326 5958
rect 8350 5956 8406 5958
rect 8430 5956 8486 5958
rect 8510 5956 8566 5958
rect 8206 5616 8262 5672
rect 8850 5208 8906 5264
rect 8270 4922 8326 4924
rect 8350 4922 8406 4924
rect 8430 4922 8486 4924
rect 8510 4922 8566 4924
rect 8270 4870 8296 4922
rect 8296 4870 8326 4922
rect 8350 4870 8360 4922
rect 8360 4870 8406 4922
rect 8430 4870 8476 4922
rect 8476 4870 8486 4922
rect 8510 4870 8540 4922
rect 8540 4870 8566 4922
rect 8270 4868 8326 4870
rect 8350 4868 8406 4870
rect 8430 4868 8486 4870
rect 8510 4868 8566 4870
rect 8666 4528 8722 4584
rect 8270 3834 8326 3836
rect 8350 3834 8406 3836
rect 8430 3834 8486 3836
rect 8510 3834 8566 3836
rect 8270 3782 8296 3834
rect 8296 3782 8326 3834
rect 8350 3782 8360 3834
rect 8360 3782 8406 3834
rect 8430 3782 8476 3834
rect 8476 3782 8486 3834
rect 8510 3782 8540 3834
rect 8540 3782 8566 3834
rect 8270 3780 8326 3782
rect 8350 3780 8406 3782
rect 8430 3780 8486 3782
rect 8510 3780 8566 3782
rect 7010 3476 7012 3496
rect 7012 3476 7064 3496
rect 7064 3476 7066 3496
rect 7010 3440 7066 3476
rect 7102 2916 7158 2952
rect 7102 2896 7104 2916
rect 7104 2896 7156 2916
rect 7156 2896 7158 2916
rect 8114 3476 8116 3496
rect 8116 3476 8168 3496
rect 8168 3476 8170 3496
rect 8114 3440 8170 3476
rect 10708 15258 10764 15260
rect 10788 15258 10844 15260
rect 10868 15258 10924 15260
rect 10948 15258 11004 15260
rect 10708 15206 10734 15258
rect 10734 15206 10764 15258
rect 10788 15206 10798 15258
rect 10798 15206 10844 15258
rect 10868 15206 10914 15258
rect 10914 15206 10924 15258
rect 10948 15206 10978 15258
rect 10978 15206 11004 15258
rect 10708 15204 10764 15206
rect 10788 15204 10844 15206
rect 10868 15204 10924 15206
rect 10948 15204 11004 15206
rect 10708 14170 10764 14172
rect 10788 14170 10844 14172
rect 10868 14170 10924 14172
rect 10948 14170 11004 14172
rect 10708 14118 10734 14170
rect 10734 14118 10764 14170
rect 10788 14118 10798 14170
rect 10798 14118 10844 14170
rect 10868 14118 10914 14170
rect 10914 14118 10924 14170
rect 10948 14118 10978 14170
rect 10978 14118 11004 14170
rect 10708 14116 10764 14118
rect 10788 14116 10844 14118
rect 10868 14116 10924 14118
rect 10948 14116 11004 14118
rect 13146 15802 13202 15804
rect 13226 15802 13282 15804
rect 13306 15802 13362 15804
rect 13386 15802 13442 15804
rect 13146 15750 13172 15802
rect 13172 15750 13202 15802
rect 13226 15750 13236 15802
rect 13236 15750 13282 15802
rect 13306 15750 13352 15802
rect 13352 15750 13362 15802
rect 13386 15750 13416 15802
rect 13416 15750 13442 15802
rect 13146 15748 13202 15750
rect 13226 15748 13282 15750
rect 13306 15748 13362 15750
rect 13386 15748 13442 15750
rect 9402 9424 9458 9480
rect 9678 9460 9680 9480
rect 9680 9460 9732 9480
rect 9732 9460 9734 9480
rect 9678 9424 9734 9460
rect 9126 6024 9182 6080
rect 9586 6568 9642 6624
rect 9586 6452 9642 6488
rect 9586 6432 9588 6452
rect 9588 6432 9640 6452
rect 9640 6432 9642 6452
rect 9310 6332 9312 6352
rect 9312 6332 9364 6352
rect 9364 6332 9366 6352
rect 9310 6296 9366 6332
rect 10708 13082 10764 13084
rect 10788 13082 10844 13084
rect 10868 13082 10924 13084
rect 10948 13082 11004 13084
rect 10708 13030 10734 13082
rect 10734 13030 10764 13082
rect 10788 13030 10798 13082
rect 10798 13030 10844 13082
rect 10868 13030 10914 13082
rect 10914 13030 10924 13082
rect 10948 13030 10978 13082
rect 10978 13030 11004 13082
rect 10708 13028 10764 13030
rect 10788 13028 10844 13030
rect 10868 13028 10924 13030
rect 10948 13028 11004 13030
rect 10708 11994 10764 11996
rect 10788 11994 10844 11996
rect 10868 11994 10924 11996
rect 10948 11994 11004 11996
rect 10708 11942 10734 11994
rect 10734 11942 10764 11994
rect 10788 11942 10798 11994
rect 10798 11942 10844 11994
rect 10868 11942 10914 11994
rect 10914 11942 10924 11994
rect 10948 11942 10978 11994
rect 10978 11942 11004 11994
rect 10708 11940 10764 11942
rect 10788 11940 10844 11942
rect 10868 11940 10924 11942
rect 10948 11940 11004 11942
rect 9586 6196 9588 6216
rect 9588 6196 9640 6216
rect 9640 6196 9642 6216
rect 9586 6160 9642 6196
rect 9494 6024 9550 6080
rect 9770 5636 9826 5672
rect 9770 5616 9772 5636
rect 9772 5616 9824 5636
rect 9824 5616 9826 5636
rect 9770 5072 9826 5128
rect 9678 4392 9734 4448
rect 8270 2746 8326 2748
rect 8350 2746 8406 2748
rect 8430 2746 8486 2748
rect 8510 2746 8566 2748
rect 8270 2694 8296 2746
rect 8296 2694 8326 2746
rect 8350 2694 8360 2746
rect 8360 2694 8406 2746
rect 8430 2694 8476 2746
rect 8476 2694 8486 2746
rect 8510 2694 8540 2746
rect 8540 2694 8566 2746
rect 8270 2692 8326 2694
rect 8350 2692 8406 2694
rect 8430 2692 8486 2694
rect 8510 2692 8566 2694
rect 10708 10906 10764 10908
rect 10788 10906 10844 10908
rect 10868 10906 10924 10908
rect 10948 10906 11004 10908
rect 10708 10854 10734 10906
rect 10734 10854 10764 10906
rect 10788 10854 10798 10906
rect 10798 10854 10844 10906
rect 10868 10854 10914 10906
rect 10914 10854 10924 10906
rect 10948 10854 10978 10906
rect 10978 10854 11004 10906
rect 10708 10852 10764 10854
rect 10788 10852 10844 10854
rect 10868 10852 10924 10854
rect 10948 10852 11004 10854
rect 10708 9818 10764 9820
rect 10788 9818 10844 9820
rect 10868 9818 10924 9820
rect 10948 9818 11004 9820
rect 10708 9766 10734 9818
rect 10734 9766 10764 9818
rect 10788 9766 10798 9818
rect 10798 9766 10844 9818
rect 10868 9766 10914 9818
rect 10914 9766 10924 9818
rect 10948 9766 10978 9818
rect 10978 9766 11004 9818
rect 10708 9764 10764 9766
rect 10788 9764 10844 9766
rect 10868 9764 10924 9766
rect 10948 9764 11004 9766
rect 11150 9560 11206 9616
rect 10708 8730 10764 8732
rect 10788 8730 10844 8732
rect 10868 8730 10924 8732
rect 10948 8730 11004 8732
rect 10708 8678 10734 8730
rect 10734 8678 10764 8730
rect 10788 8678 10798 8730
rect 10798 8678 10844 8730
rect 10868 8678 10914 8730
rect 10914 8678 10924 8730
rect 10948 8678 10978 8730
rect 10978 8678 11004 8730
rect 10708 8676 10764 8678
rect 10788 8676 10844 8678
rect 10868 8676 10924 8678
rect 10948 8676 11004 8678
rect 10506 8084 10562 8120
rect 10506 8064 10508 8084
rect 10508 8064 10560 8084
rect 10560 8064 10562 8084
rect 10708 7642 10764 7644
rect 10788 7642 10844 7644
rect 10868 7642 10924 7644
rect 10948 7642 11004 7644
rect 10708 7590 10734 7642
rect 10734 7590 10764 7642
rect 10788 7590 10798 7642
rect 10798 7590 10844 7642
rect 10868 7590 10914 7642
rect 10914 7590 10924 7642
rect 10948 7590 10978 7642
rect 10978 7590 11004 7642
rect 10708 7588 10764 7590
rect 10788 7588 10844 7590
rect 10868 7588 10924 7590
rect 10948 7588 11004 7590
rect 10708 6554 10764 6556
rect 10788 6554 10844 6556
rect 10868 6554 10924 6556
rect 10948 6554 11004 6556
rect 10708 6502 10734 6554
rect 10734 6502 10764 6554
rect 10788 6502 10798 6554
rect 10798 6502 10844 6554
rect 10868 6502 10914 6554
rect 10914 6502 10924 6554
rect 10948 6502 10978 6554
rect 10978 6502 11004 6554
rect 10708 6500 10764 6502
rect 10788 6500 10844 6502
rect 10868 6500 10924 6502
rect 10948 6500 11004 6502
rect 10966 5752 11022 5808
rect 10708 5466 10764 5468
rect 10788 5466 10844 5468
rect 10868 5466 10924 5468
rect 10948 5466 11004 5468
rect 10708 5414 10734 5466
rect 10734 5414 10764 5466
rect 10788 5414 10798 5466
rect 10798 5414 10844 5466
rect 10868 5414 10914 5466
rect 10914 5414 10924 5466
rect 10948 5414 10978 5466
rect 10978 5414 11004 5466
rect 10708 5412 10764 5414
rect 10788 5412 10844 5414
rect 10868 5412 10924 5414
rect 10948 5412 11004 5414
rect 10598 4936 10654 4992
rect 11610 9424 11666 9480
rect 12162 10004 12164 10024
rect 12164 10004 12216 10024
rect 12216 10004 12218 10024
rect 12162 9968 12218 10004
rect 13146 14714 13202 14716
rect 13226 14714 13282 14716
rect 13306 14714 13362 14716
rect 13386 14714 13442 14716
rect 13146 14662 13172 14714
rect 13172 14662 13202 14714
rect 13226 14662 13236 14714
rect 13236 14662 13282 14714
rect 13306 14662 13352 14714
rect 13352 14662 13362 14714
rect 13386 14662 13416 14714
rect 13416 14662 13442 14714
rect 13146 14660 13202 14662
rect 13226 14660 13282 14662
rect 13306 14660 13362 14662
rect 13386 14660 13442 14662
rect 13146 13626 13202 13628
rect 13226 13626 13282 13628
rect 13306 13626 13362 13628
rect 13386 13626 13442 13628
rect 13146 13574 13172 13626
rect 13172 13574 13202 13626
rect 13226 13574 13236 13626
rect 13236 13574 13282 13626
rect 13306 13574 13352 13626
rect 13352 13574 13362 13626
rect 13386 13574 13416 13626
rect 13416 13574 13442 13626
rect 13146 13572 13202 13574
rect 13226 13572 13282 13574
rect 13306 13572 13362 13574
rect 13386 13572 13442 13574
rect 13146 12538 13202 12540
rect 13226 12538 13282 12540
rect 13306 12538 13362 12540
rect 13386 12538 13442 12540
rect 13146 12486 13172 12538
rect 13172 12486 13202 12538
rect 13226 12486 13236 12538
rect 13236 12486 13282 12538
rect 13306 12486 13352 12538
rect 13352 12486 13362 12538
rect 13386 12486 13416 12538
rect 13416 12486 13442 12538
rect 13146 12484 13202 12486
rect 13226 12484 13282 12486
rect 13306 12484 13362 12486
rect 13386 12484 13442 12486
rect 13146 11450 13202 11452
rect 13226 11450 13282 11452
rect 13306 11450 13362 11452
rect 13386 11450 13442 11452
rect 13146 11398 13172 11450
rect 13172 11398 13202 11450
rect 13226 11398 13236 11450
rect 13236 11398 13282 11450
rect 13306 11398 13352 11450
rect 13352 11398 13362 11450
rect 13386 11398 13416 11450
rect 13416 11398 13442 11450
rect 13146 11396 13202 11398
rect 13226 11396 13282 11398
rect 13306 11396 13362 11398
rect 13386 11396 13442 11398
rect 12438 10140 12440 10160
rect 12440 10140 12492 10160
rect 12492 10140 12494 10160
rect 12438 10104 12494 10140
rect 11518 5244 11520 5264
rect 11520 5244 11572 5264
rect 11572 5244 11574 5264
rect 11518 5208 11574 5244
rect 11610 5072 11666 5128
rect 11426 4528 11482 4584
rect 10708 4378 10764 4380
rect 10788 4378 10844 4380
rect 10868 4378 10924 4380
rect 10948 4378 11004 4380
rect 10708 4326 10734 4378
rect 10734 4326 10764 4378
rect 10788 4326 10798 4378
rect 10798 4326 10844 4378
rect 10868 4326 10914 4378
rect 10914 4326 10924 4378
rect 10948 4326 10978 4378
rect 10978 4326 11004 4378
rect 10708 4324 10764 4326
rect 10788 4324 10844 4326
rect 10868 4324 10924 4326
rect 10948 4324 11004 4326
rect 12438 7928 12494 7984
rect 12070 5752 12126 5808
rect 11978 5072 12034 5128
rect 12438 5228 12494 5264
rect 12438 5208 12440 5228
rect 12440 5208 12492 5228
rect 12492 5208 12494 5228
rect 10708 3290 10764 3292
rect 10788 3290 10844 3292
rect 10868 3290 10924 3292
rect 10948 3290 11004 3292
rect 10708 3238 10734 3290
rect 10734 3238 10764 3290
rect 10788 3238 10798 3290
rect 10798 3238 10844 3290
rect 10868 3238 10914 3290
rect 10914 3238 10924 3290
rect 10948 3238 10978 3290
rect 10978 3238 11004 3290
rect 10708 3236 10764 3238
rect 10788 3236 10844 3238
rect 10868 3236 10924 3238
rect 10948 3236 11004 3238
rect 12162 2896 12218 2952
rect 13146 10362 13202 10364
rect 13226 10362 13282 10364
rect 13306 10362 13362 10364
rect 13386 10362 13442 10364
rect 13146 10310 13172 10362
rect 13172 10310 13202 10362
rect 13226 10310 13236 10362
rect 13236 10310 13282 10362
rect 13306 10310 13352 10362
rect 13352 10310 13362 10362
rect 13386 10310 13416 10362
rect 13416 10310 13442 10362
rect 13146 10308 13202 10310
rect 13226 10308 13282 10310
rect 13306 10308 13362 10310
rect 13386 10308 13442 10310
rect 13082 10140 13084 10160
rect 13084 10140 13136 10160
rect 13136 10140 13138 10160
rect 13082 10104 13138 10140
rect 13358 9988 13414 10024
rect 13358 9968 13360 9988
rect 13360 9968 13412 9988
rect 13412 9968 13414 9988
rect 13146 9274 13202 9276
rect 13226 9274 13282 9276
rect 13306 9274 13362 9276
rect 13386 9274 13442 9276
rect 13146 9222 13172 9274
rect 13172 9222 13202 9274
rect 13226 9222 13236 9274
rect 13236 9222 13282 9274
rect 13306 9222 13352 9274
rect 13352 9222 13362 9274
rect 13386 9222 13416 9274
rect 13416 9222 13442 9274
rect 13146 9220 13202 9222
rect 13226 9220 13282 9222
rect 13306 9220 13362 9222
rect 13386 9220 13442 9222
rect 12806 8064 12862 8120
rect 13146 8186 13202 8188
rect 13226 8186 13282 8188
rect 13306 8186 13362 8188
rect 13386 8186 13442 8188
rect 13146 8134 13172 8186
rect 13172 8134 13202 8186
rect 13226 8134 13236 8186
rect 13236 8134 13282 8186
rect 13306 8134 13352 8186
rect 13352 8134 13362 8186
rect 13386 8134 13416 8186
rect 13416 8134 13442 8186
rect 13146 8132 13202 8134
rect 13226 8132 13282 8134
rect 13306 8132 13362 8134
rect 13386 8132 13442 8134
rect 13146 7098 13202 7100
rect 13226 7098 13282 7100
rect 13306 7098 13362 7100
rect 13386 7098 13442 7100
rect 13146 7046 13172 7098
rect 13172 7046 13202 7098
rect 13226 7046 13236 7098
rect 13236 7046 13282 7098
rect 13306 7046 13352 7098
rect 13352 7046 13362 7098
rect 13386 7046 13416 7098
rect 13416 7046 13442 7098
rect 13146 7044 13202 7046
rect 13226 7044 13282 7046
rect 13306 7044 13362 7046
rect 13386 7044 13442 7046
rect 12806 5752 12862 5808
rect 13146 6010 13202 6012
rect 13226 6010 13282 6012
rect 13306 6010 13362 6012
rect 13386 6010 13442 6012
rect 13146 5958 13172 6010
rect 13172 5958 13202 6010
rect 13226 5958 13236 6010
rect 13236 5958 13282 6010
rect 13306 5958 13352 6010
rect 13352 5958 13362 6010
rect 13386 5958 13416 6010
rect 13416 5958 13442 6010
rect 13146 5956 13202 5958
rect 13226 5956 13282 5958
rect 13306 5956 13362 5958
rect 13386 5956 13442 5958
rect 13146 4922 13202 4924
rect 13226 4922 13282 4924
rect 13306 4922 13362 4924
rect 13386 4922 13442 4924
rect 13146 4870 13172 4922
rect 13172 4870 13202 4922
rect 13226 4870 13236 4922
rect 13236 4870 13282 4922
rect 13306 4870 13352 4922
rect 13352 4870 13362 4922
rect 13386 4870 13416 4922
rect 13416 4870 13442 4922
rect 13146 4868 13202 4870
rect 13226 4868 13282 4870
rect 13306 4868 13362 4870
rect 13386 4868 13442 4870
rect 12898 4664 12954 4720
rect 13266 4664 13322 4720
rect 13910 5616 13966 5672
rect 13146 3834 13202 3836
rect 13226 3834 13282 3836
rect 13306 3834 13362 3836
rect 13386 3834 13442 3836
rect 13146 3782 13172 3834
rect 13172 3782 13202 3834
rect 13226 3782 13236 3834
rect 13236 3782 13282 3834
rect 13306 3782 13352 3834
rect 13352 3782 13362 3834
rect 13386 3782 13416 3834
rect 13416 3782 13442 3834
rect 13146 3780 13202 3782
rect 13226 3780 13282 3782
rect 13306 3780 13362 3782
rect 13386 3780 13442 3782
rect 13146 2746 13202 2748
rect 13226 2746 13282 2748
rect 13306 2746 13362 2748
rect 13386 2746 13442 2748
rect 13146 2694 13172 2746
rect 13172 2694 13202 2746
rect 13226 2694 13236 2746
rect 13236 2694 13282 2746
rect 13306 2694 13352 2746
rect 13352 2694 13362 2746
rect 13386 2694 13416 2746
rect 13416 2694 13442 2746
rect 13146 2692 13202 2694
rect 13226 2692 13282 2694
rect 13306 2692 13362 2694
rect 13386 2692 13442 2694
rect 13542 2488 13598 2544
rect 15014 16108 15070 16144
rect 15014 16088 15016 16108
rect 15016 16088 15068 16108
rect 15068 16088 15070 16108
rect 15014 13368 15070 13424
rect 14462 4528 14518 4584
rect 14922 10648 14978 10704
rect 15014 5228 15070 5264
rect 15014 5208 15016 5228
rect 15016 5208 15068 5228
rect 15068 5208 15070 5228
rect 10708 2202 10764 2204
rect 10788 2202 10844 2204
rect 10868 2202 10924 2204
rect 10948 2202 11004 2204
rect 10708 2150 10734 2202
rect 10734 2150 10764 2202
rect 10788 2150 10798 2202
rect 10798 2150 10844 2202
rect 10868 2150 10914 2202
rect 10914 2150 10924 2202
rect 10948 2150 10978 2202
rect 10978 2150 11004 2202
rect 10708 2148 10764 2150
rect 10788 2148 10844 2150
rect 10868 2148 10924 2150
rect 10948 2148 11004 2150
<< metal3 >>
rect 0 16418 800 16448
rect 1393 16418 1459 16421
rect 0 16416 1459 16418
rect 0 16360 1398 16416
rect 1454 16360 1459 16416
rect 0 16358 1459 16360
rect 0 16328 800 16358
rect 1393 16355 1459 16358
rect 5820 16352 6140 16353
rect 5820 16288 5828 16352
rect 5892 16288 5908 16352
rect 5972 16288 5988 16352
rect 6052 16288 6068 16352
rect 6132 16288 6140 16352
rect 5820 16287 6140 16288
rect 10696 16352 11016 16353
rect 10696 16288 10704 16352
rect 10768 16288 10784 16352
rect 10848 16288 10864 16352
rect 10928 16288 10944 16352
rect 11008 16288 11016 16352
rect 10696 16287 11016 16288
rect 15009 16146 15075 16149
rect 16071 16146 16871 16176
rect 15009 16144 16871 16146
rect 15009 16088 15014 16144
rect 15070 16088 16871 16144
rect 15009 16086 16871 16088
rect 15009 16083 15075 16086
rect 16071 16056 16871 16086
rect 3382 15808 3702 15809
rect 3382 15744 3390 15808
rect 3454 15744 3470 15808
rect 3534 15744 3550 15808
rect 3614 15744 3630 15808
rect 3694 15744 3702 15808
rect 3382 15743 3702 15744
rect 8258 15808 8578 15809
rect 8258 15744 8266 15808
rect 8330 15744 8346 15808
rect 8410 15744 8426 15808
rect 8490 15744 8506 15808
rect 8570 15744 8578 15808
rect 8258 15743 8578 15744
rect 13134 15808 13454 15809
rect 13134 15744 13142 15808
rect 13206 15744 13222 15808
rect 13286 15744 13302 15808
rect 13366 15744 13382 15808
rect 13446 15744 13454 15808
rect 13134 15743 13454 15744
rect 5820 15264 6140 15265
rect 5820 15200 5828 15264
rect 5892 15200 5908 15264
rect 5972 15200 5988 15264
rect 6052 15200 6068 15264
rect 6132 15200 6140 15264
rect 5820 15199 6140 15200
rect 10696 15264 11016 15265
rect 10696 15200 10704 15264
rect 10768 15200 10784 15264
rect 10848 15200 10864 15264
rect 10928 15200 10944 15264
rect 11008 15200 11016 15264
rect 10696 15199 11016 15200
rect 3382 14720 3702 14721
rect 3382 14656 3390 14720
rect 3454 14656 3470 14720
rect 3534 14656 3550 14720
rect 3614 14656 3630 14720
rect 3694 14656 3702 14720
rect 3382 14655 3702 14656
rect 8258 14720 8578 14721
rect 8258 14656 8266 14720
rect 8330 14656 8346 14720
rect 8410 14656 8426 14720
rect 8490 14656 8506 14720
rect 8570 14656 8578 14720
rect 8258 14655 8578 14656
rect 13134 14720 13454 14721
rect 13134 14656 13142 14720
rect 13206 14656 13222 14720
rect 13286 14656 13302 14720
rect 13366 14656 13382 14720
rect 13446 14656 13454 14720
rect 13134 14655 13454 14656
rect 5820 14176 6140 14177
rect 5820 14112 5828 14176
rect 5892 14112 5908 14176
rect 5972 14112 5988 14176
rect 6052 14112 6068 14176
rect 6132 14112 6140 14176
rect 5820 14111 6140 14112
rect 10696 14176 11016 14177
rect 10696 14112 10704 14176
rect 10768 14112 10784 14176
rect 10848 14112 10864 14176
rect 10928 14112 10944 14176
rect 11008 14112 11016 14176
rect 10696 14111 11016 14112
rect 0 13698 800 13728
rect 1853 13698 1919 13701
rect 0 13696 1919 13698
rect 0 13640 1858 13696
rect 1914 13640 1919 13696
rect 0 13638 1919 13640
rect 0 13608 800 13638
rect 1853 13635 1919 13638
rect 3382 13632 3702 13633
rect 3382 13568 3390 13632
rect 3454 13568 3470 13632
rect 3534 13568 3550 13632
rect 3614 13568 3630 13632
rect 3694 13568 3702 13632
rect 3382 13567 3702 13568
rect 8258 13632 8578 13633
rect 8258 13568 8266 13632
rect 8330 13568 8346 13632
rect 8410 13568 8426 13632
rect 8490 13568 8506 13632
rect 8570 13568 8578 13632
rect 8258 13567 8578 13568
rect 13134 13632 13454 13633
rect 13134 13568 13142 13632
rect 13206 13568 13222 13632
rect 13286 13568 13302 13632
rect 13366 13568 13382 13632
rect 13446 13568 13454 13632
rect 13134 13567 13454 13568
rect 15009 13426 15075 13429
rect 16071 13426 16871 13456
rect 15009 13424 16871 13426
rect 15009 13368 15014 13424
rect 15070 13368 16871 13424
rect 15009 13366 16871 13368
rect 15009 13363 15075 13366
rect 16071 13336 16871 13366
rect 5820 13088 6140 13089
rect 5820 13024 5828 13088
rect 5892 13024 5908 13088
rect 5972 13024 5988 13088
rect 6052 13024 6068 13088
rect 6132 13024 6140 13088
rect 5820 13023 6140 13024
rect 10696 13088 11016 13089
rect 10696 13024 10704 13088
rect 10768 13024 10784 13088
rect 10848 13024 10864 13088
rect 10928 13024 10944 13088
rect 11008 13024 11016 13088
rect 10696 13023 11016 13024
rect 3382 12544 3702 12545
rect 3382 12480 3390 12544
rect 3454 12480 3470 12544
rect 3534 12480 3550 12544
rect 3614 12480 3630 12544
rect 3694 12480 3702 12544
rect 3382 12479 3702 12480
rect 8258 12544 8578 12545
rect 8258 12480 8266 12544
rect 8330 12480 8346 12544
rect 8410 12480 8426 12544
rect 8490 12480 8506 12544
rect 8570 12480 8578 12544
rect 8258 12479 8578 12480
rect 13134 12544 13454 12545
rect 13134 12480 13142 12544
rect 13206 12480 13222 12544
rect 13286 12480 13302 12544
rect 13366 12480 13382 12544
rect 13446 12480 13454 12544
rect 13134 12479 13454 12480
rect 5820 12000 6140 12001
rect 5820 11936 5828 12000
rect 5892 11936 5908 12000
rect 5972 11936 5988 12000
rect 6052 11936 6068 12000
rect 6132 11936 6140 12000
rect 5820 11935 6140 11936
rect 10696 12000 11016 12001
rect 10696 11936 10704 12000
rect 10768 11936 10784 12000
rect 10848 11936 10864 12000
rect 10928 11936 10944 12000
rect 11008 11936 11016 12000
rect 10696 11935 11016 11936
rect 3382 11456 3702 11457
rect 3382 11392 3390 11456
rect 3454 11392 3470 11456
rect 3534 11392 3550 11456
rect 3614 11392 3630 11456
rect 3694 11392 3702 11456
rect 3382 11391 3702 11392
rect 8258 11456 8578 11457
rect 8258 11392 8266 11456
rect 8330 11392 8346 11456
rect 8410 11392 8426 11456
rect 8490 11392 8506 11456
rect 8570 11392 8578 11456
rect 8258 11391 8578 11392
rect 13134 11456 13454 11457
rect 13134 11392 13142 11456
rect 13206 11392 13222 11456
rect 13286 11392 13302 11456
rect 13366 11392 13382 11456
rect 13446 11392 13454 11456
rect 13134 11391 13454 11392
rect 0 10978 800 11008
rect 1853 10978 1919 10981
rect 0 10976 1919 10978
rect 0 10920 1858 10976
rect 1914 10920 1919 10976
rect 0 10918 1919 10920
rect 0 10888 800 10918
rect 1853 10915 1919 10918
rect 5820 10912 6140 10913
rect 5820 10848 5828 10912
rect 5892 10848 5908 10912
rect 5972 10848 5988 10912
rect 6052 10848 6068 10912
rect 6132 10848 6140 10912
rect 5820 10847 6140 10848
rect 10696 10912 11016 10913
rect 10696 10848 10704 10912
rect 10768 10848 10784 10912
rect 10848 10848 10864 10912
rect 10928 10848 10944 10912
rect 11008 10848 11016 10912
rect 10696 10847 11016 10848
rect 5717 10706 5783 10709
rect 7189 10706 7255 10709
rect 5717 10704 7255 10706
rect 5717 10648 5722 10704
rect 5778 10648 7194 10704
rect 7250 10648 7255 10704
rect 5717 10646 7255 10648
rect 5717 10643 5783 10646
rect 7189 10643 7255 10646
rect 14917 10706 14983 10709
rect 16071 10706 16871 10736
rect 14917 10704 16871 10706
rect 14917 10648 14922 10704
rect 14978 10648 16871 10704
rect 14917 10646 16871 10648
rect 14917 10643 14983 10646
rect 16071 10616 16871 10646
rect 3382 10368 3702 10369
rect 3382 10304 3390 10368
rect 3454 10304 3470 10368
rect 3534 10304 3550 10368
rect 3614 10304 3630 10368
rect 3694 10304 3702 10368
rect 3382 10303 3702 10304
rect 8258 10368 8578 10369
rect 8258 10304 8266 10368
rect 8330 10304 8346 10368
rect 8410 10304 8426 10368
rect 8490 10304 8506 10368
rect 8570 10304 8578 10368
rect 8258 10303 8578 10304
rect 13134 10368 13454 10369
rect 13134 10304 13142 10368
rect 13206 10304 13222 10368
rect 13286 10304 13302 10368
rect 13366 10304 13382 10368
rect 13446 10304 13454 10368
rect 13134 10303 13454 10304
rect 12433 10162 12499 10165
rect 13077 10162 13143 10165
rect 12433 10160 13143 10162
rect 12433 10104 12438 10160
rect 12494 10104 13082 10160
rect 13138 10104 13143 10160
rect 12433 10102 13143 10104
rect 12433 10099 12499 10102
rect 13077 10099 13143 10102
rect 12157 10026 12223 10029
rect 13353 10026 13419 10029
rect 12157 10024 13419 10026
rect 12157 9968 12162 10024
rect 12218 9968 13358 10024
rect 13414 9968 13419 10024
rect 12157 9966 13419 9968
rect 12157 9963 12223 9966
rect 13353 9963 13419 9966
rect 5820 9824 6140 9825
rect 5820 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6140 9824
rect 5820 9759 6140 9760
rect 10696 9824 11016 9825
rect 10696 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11016 9824
rect 10696 9759 11016 9760
rect 5625 9618 5691 9621
rect 11145 9618 11211 9621
rect 5625 9616 11211 9618
rect 5625 9560 5630 9616
rect 5686 9560 11150 9616
rect 11206 9560 11211 9616
rect 5625 9558 11211 9560
rect 5625 9555 5691 9558
rect 11145 9555 11211 9558
rect 3785 9482 3851 9485
rect 5717 9482 5783 9485
rect 3785 9480 5783 9482
rect 3785 9424 3790 9480
rect 3846 9424 5722 9480
rect 5778 9424 5783 9480
rect 3785 9422 5783 9424
rect 3785 9419 3851 9422
rect 5717 9419 5783 9422
rect 8109 9482 8175 9485
rect 9397 9482 9463 9485
rect 8109 9480 9463 9482
rect 8109 9424 8114 9480
rect 8170 9424 9402 9480
rect 9458 9424 9463 9480
rect 8109 9422 9463 9424
rect 8109 9419 8175 9422
rect 9397 9419 9463 9422
rect 9673 9482 9739 9485
rect 11605 9482 11671 9485
rect 9673 9480 11671 9482
rect 9673 9424 9678 9480
rect 9734 9424 11610 9480
rect 11666 9424 11671 9480
rect 9673 9422 11671 9424
rect 9673 9419 9739 9422
rect 11605 9419 11671 9422
rect 3382 9280 3702 9281
rect 3382 9216 3390 9280
rect 3454 9216 3470 9280
rect 3534 9216 3550 9280
rect 3614 9216 3630 9280
rect 3694 9216 3702 9280
rect 3382 9215 3702 9216
rect 8258 9280 8578 9281
rect 8258 9216 8266 9280
rect 8330 9216 8346 9280
rect 8410 9216 8426 9280
rect 8490 9216 8506 9280
rect 8570 9216 8578 9280
rect 8258 9215 8578 9216
rect 13134 9280 13454 9281
rect 13134 9216 13142 9280
rect 13206 9216 13222 9280
rect 13286 9216 13302 9280
rect 13366 9216 13382 9280
rect 13446 9216 13454 9280
rect 13134 9215 13454 9216
rect 5820 8736 6140 8737
rect 5820 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6140 8736
rect 5820 8671 6140 8672
rect 10696 8736 11016 8737
rect 10696 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11016 8736
rect 10696 8671 11016 8672
rect 0 8258 800 8288
rect 2865 8258 2931 8261
rect 0 8256 2931 8258
rect 0 8200 2870 8256
rect 2926 8200 2931 8256
rect 0 8198 2931 8200
rect 0 8168 800 8198
rect 2865 8195 2931 8198
rect 3382 8192 3702 8193
rect 3382 8128 3390 8192
rect 3454 8128 3470 8192
rect 3534 8128 3550 8192
rect 3614 8128 3630 8192
rect 3694 8128 3702 8192
rect 3382 8127 3702 8128
rect 8258 8192 8578 8193
rect 8258 8128 8266 8192
rect 8330 8128 8346 8192
rect 8410 8128 8426 8192
rect 8490 8128 8506 8192
rect 8570 8128 8578 8192
rect 8258 8127 8578 8128
rect 13134 8192 13454 8193
rect 13134 8128 13142 8192
rect 13206 8128 13222 8192
rect 13286 8128 13302 8192
rect 13366 8128 13382 8192
rect 13446 8128 13454 8192
rect 13134 8127 13454 8128
rect 10501 8122 10567 8125
rect 12801 8122 12867 8125
rect 10501 8120 12867 8122
rect 10501 8064 10506 8120
rect 10562 8064 12806 8120
rect 12862 8064 12867 8120
rect 10501 8062 12867 8064
rect 10501 8059 10567 8062
rect 12801 8059 12867 8062
rect 12433 7986 12499 7989
rect 16071 7986 16871 8016
rect 12433 7984 16871 7986
rect 12433 7928 12438 7984
rect 12494 7928 16871 7984
rect 12433 7926 16871 7928
rect 12433 7923 12499 7926
rect 16071 7896 16871 7926
rect 5820 7648 6140 7649
rect 5820 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6140 7648
rect 5820 7583 6140 7584
rect 10696 7648 11016 7649
rect 10696 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11016 7648
rect 10696 7583 11016 7584
rect 3382 7104 3702 7105
rect 3382 7040 3390 7104
rect 3454 7040 3470 7104
rect 3534 7040 3550 7104
rect 3614 7040 3630 7104
rect 3694 7040 3702 7104
rect 3382 7039 3702 7040
rect 8258 7104 8578 7105
rect 8258 7040 8266 7104
rect 8330 7040 8346 7104
rect 8410 7040 8426 7104
rect 8490 7040 8506 7104
rect 8570 7040 8578 7104
rect 8258 7039 8578 7040
rect 13134 7104 13454 7105
rect 13134 7040 13142 7104
rect 13206 7040 13222 7104
rect 13286 7040 13302 7104
rect 13366 7040 13382 7104
rect 13446 7040 13454 7104
rect 13134 7039 13454 7040
rect 8569 6626 8635 6629
rect 9581 6626 9647 6629
rect 8569 6624 9647 6626
rect 8569 6568 8574 6624
rect 8630 6568 9586 6624
rect 9642 6568 9647 6624
rect 8569 6566 9647 6568
rect 8569 6563 8635 6566
rect 9581 6563 9647 6566
rect 5820 6560 6140 6561
rect 5820 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6140 6560
rect 5820 6495 6140 6496
rect 10696 6560 11016 6561
rect 10696 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11016 6560
rect 10696 6495 11016 6496
rect 7097 6490 7163 6493
rect 9581 6490 9647 6493
rect 7097 6488 9647 6490
rect 7097 6432 7102 6488
rect 7158 6432 9586 6488
rect 9642 6432 9647 6488
rect 7097 6430 9647 6432
rect 7097 6427 7163 6430
rect 9581 6427 9647 6430
rect 7189 6354 7255 6357
rect 9305 6354 9371 6357
rect 7189 6352 9371 6354
rect 7189 6296 7194 6352
rect 7250 6296 9310 6352
rect 9366 6296 9371 6352
rect 7189 6294 9371 6296
rect 7189 6291 7255 6294
rect 9305 6291 9371 6294
rect 8385 6218 8451 6221
rect 9581 6218 9647 6221
rect 8385 6216 9647 6218
rect 8385 6160 8390 6216
rect 8446 6160 9586 6216
rect 9642 6160 9647 6216
rect 8385 6158 9647 6160
rect 8385 6155 8451 6158
rect 9581 6155 9647 6158
rect 9121 6082 9187 6085
rect 9489 6082 9555 6085
rect 9121 6080 9555 6082
rect 9121 6024 9126 6080
rect 9182 6024 9494 6080
rect 9550 6024 9555 6080
rect 9121 6022 9555 6024
rect 9121 6019 9187 6022
rect 9489 6019 9555 6022
rect 3382 6016 3702 6017
rect 3382 5952 3390 6016
rect 3454 5952 3470 6016
rect 3534 5952 3550 6016
rect 3614 5952 3630 6016
rect 3694 5952 3702 6016
rect 3382 5951 3702 5952
rect 8258 6016 8578 6017
rect 8258 5952 8266 6016
rect 8330 5952 8346 6016
rect 8410 5952 8426 6016
rect 8490 5952 8506 6016
rect 8570 5952 8578 6016
rect 8258 5951 8578 5952
rect 13134 6016 13454 6017
rect 13134 5952 13142 6016
rect 13206 5952 13222 6016
rect 13286 5952 13302 6016
rect 13366 5952 13382 6016
rect 13446 5952 13454 6016
rect 13134 5951 13454 5952
rect 10961 5810 11027 5813
rect 12065 5810 12131 5813
rect 12801 5810 12867 5813
rect 10961 5808 12867 5810
rect 10961 5752 10966 5808
rect 11022 5752 12070 5808
rect 12126 5752 12806 5808
rect 12862 5752 12867 5808
rect 10961 5750 12867 5752
rect 10961 5747 11027 5750
rect 12065 5747 12131 5750
rect 12801 5747 12867 5750
rect 2405 5674 2471 5677
rect 8201 5674 8267 5677
rect 2405 5672 8267 5674
rect 2405 5616 2410 5672
rect 2466 5616 8206 5672
rect 8262 5616 8267 5672
rect 2405 5614 8267 5616
rect 2405 5611 2471 5614
rect 8201 5611 8267 5614
rect 9765 5674 9831 5677
rect 13905 5674 13971 5677
rect 9765 5672 13971 5674
rect 9765 5616 9770 5672
rect 9826 5616 13910 5672
rect 13966 5616 13971 5672
rect 9765 5614 13971 5616
rect 9765 5611 9831 5614
rect 13905 5611 13971 5614
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 5820 5472 6140 5473
rect 5820 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6140 5472
rect 5820 5407 6140 5408
rect 10696 5472 11016 5473
rect 10696 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11016 5472
rect 10696 5407 11016 5408
rect 6177 5266 6243 5269
rect 8845 5266 8911 5269
rect 6177 5264 8911 5266
rect 6177 5208 6182 5264
rect 6238 5208 8850 5264
rect 8906 5208 8911 5264
rect 6177 5206 8911 5208
rect 6177 5203 6243 5206
rect 8845 5203 8911 5206
rect 11513 5266 11579 5269
rect 12433 5266 12499 5269
rect 11513 5264 12499 5266
rect 11513 5208 11518 5264
rect 11574 5208 12438 5264
rect 12494 5208 12499 5264
rect 11513 5206 12499 5208
rect 11513 5203 11579 5206
rect 12433 5203 12499 5206
rect 15009 5266 15075 5269
rect 16071 5266 16871 5296
rect 15009 5264 16871 5266
rect 15009 5208 15014 5264
rect 15070 5208 16871 5264
rect 15009 5206 16871 5208
rect 15009 5203 15075 5206
rect 16071 5176 16871 5206
rect 2405 5130 2471 5133
rect 9765 5130 9831 5133
rect 11605 5130 11671 5133
rect 11973 5130 12039 5133
rect 2405 5128 9690 5130
rect 2405 5072 2410 5128
rect 2466 5072 9690 5128
rect 2405 5070 9690 5072
rect 2405 5067 2471 5070
rect 9630 4994 9690 5070
rect 9765 5128 12039 5130
rect 9765 5072 9770 5128
rect 9826 5072 11610 5128
rect 11666 5072 11978 5128
rect 12034 5072 12039 5128
rect 9765 5070 12039 5072
rect 9765 5067 9831 5070
rect 11605 5067 11671 5070
rect 11973 5067 12039 5070
rect 10593 4994 10659 4997
rect 9630 4992 10659 4994
rect 9630 4936 10598 4992
rect 10654 4936 10659 4992
rect 9630 4934 10659 4936
rect 10593 4931 10659 4934
rect 3382 4928 3702 4929
rect 3382 4864 3390 4928
rect 3454 4864 3470 4928
rect 3534 4864 3550 4928
rect 3614 4864 3630 4928
rect 3694 4864 3702 4928
rect 3382 4863 3702 4864
rect 8258 4928 8578 4929
rect 8258 4864 8266 4928
rect 8330 4864 8346 4928
rect 8410 4864 8426 4928
rect 8490 4864 8506 4928
rect 8570 4864 8578 4928
rect 8258 4863 8578 4864
rect 13134 4928 13454 4929
rect 13134 4864 13142 4928
rect 13206 4864 13222 4928
rect 13286 4864 13302 4928
rect 13366 4864 13382 4928
rect 13446 4864 13454 4928
rect 13134 4863 13454 4864
rect 12893 4722 12959 4725
rect 13261 4722 13327 4725
rect 12893 4720 13327 4722
rect 12893 4664 12898 4720
rect 12954 4664 13266 4720
rect 13322 4664 13327 4720
rect 12893 4662 13327 4664
rect 12893 4659 12959 4662
rect 13261 4659 13327 4662
rect 6821 4586 6887 4589
rect 8661 4586 8727 4589
rect 6821 4584 8727 4586
rect 6821 4528 6826 4584
rect 6882 4528 8666 4584
rect 8722 4528 8727 4584
rect 6821 4526 8727 4528
rect 6821 4523 6887 4526
rect 8661 4523 8727 4526
rect 11421 4586 11487 4589
rect 14457 4586 14523 4589
rect 11421 4584 14523 4586
rect 11421 4528 11426 4584
rect 11482 4528 14462 4584
rect 14518 4528 14523 4584
rect 11421 4526 14523 4528
rect 11421 4523 11487 4526
rect 14457 4523 14523 4526
rect 6269 4450 6335 4453
rect 9673 4450 9739 4453
rect 6269 4448 9739 4450
rect 6269 4392 6274 4448
rect 6330 4392 9678 4448
rect 9734 4392 9739 4448
rect 6269 4390 9739 4392
rect 6269 4387 6335 4390
rect 9673 4387 9739 4390
rect 5820 4384 6140 4385
rect 5820 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6140 4384
rect 5820 4319 6140 4320
rect 10696 4384 11016 4385
rect 10696 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11016 4384
rect 10696 4319 11016 4320
rect 3382 3840 3702 3841
rect 3382 3776 3390 3840
rect 3454 3776 3470 3840
rect 3534 3776 3550 3840
rect 3614 3776 3630 3840
rect 3694 3776 3702 3840
rect 3382 3775 3702 3776
rect 8258 3840 8578 3841
rect 8258 3776 8266 3840
rect 8330 3776 8346 3840
rect 8410 3776 8426 3840
rect 8490 3776 8506 3840
rect 8570 3776 8578 3840
rect 8258 3775 8578 3776
rect 13134 3840 13454 3841
rect 13134 3776 13142 3840
rect 13206 3776 13222 3840
rect 13286 3776 13302 3840
rect 13366 3776 13382 3840
rect 13446 3776 13454 3840
rect 13134 3775 13454 3776
rect 7005 3498 7071 3501
rect 8109 3498 8175 3501
rect 7005 3496 8175 3498
rect 7005 3440 7010 3496
rect 7066 3440 8114 3496
rect 8170 3440 8175 3496
rect 7005 3438 8175 3440
rect 7005 3435 7071 3438
rect 8109 3435 8175 3438
rect 5820 3296 6140 3297
rect 5820 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6140 3296
rect 5820 3231 6140 3232
rect 10696 3296 11016 3297
rect 10696 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11016 3296
rect 10696 3231 11016 3232
rect 7097 2954 7163 2957
rect 12157 2954 12223 2957
rect 7097 2952 12223 2954
rect 7097 2896 7102 2952
rect 7158 2896 12162 2952
rect 12218 2896 12223 2952
rect 7097 2894 12223 2896
rect 7097 2891 7163 2894
rect 12157 2891 12223 2894
rect 0 2818 800 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 3382 2752 3702 2753
rect 3382 2688 3390 2752
rect 3454 2688 3470 2752
rect 3534 2688 3550 2752
rect 3614 2688 3630 2752
rect 3694 2688 3702 2752
rect 3382 2687 3702 2688
rect 8258 2752 8578 2753
rect 8258 2688 8266 2752
rect 8330 2688 8346 2752
rect 8410 2688 8426 2752
rect 8490 2688 8506 2752
rect 8570 2688 8578 2752
rect 8258 2687 8578 2688
rect 13134 2752 13454 2753
rect 13134 2688 13142 2752
rect 13206 2688 13222 2752
rect 13286 2688 13302 2752
rect 13366 2688 13382 2752
rect 13446 2688 13454 2752
rect 13134 2687 13454 2688
rect 13537 2546 13603 2549
rect 16071 2546 16871 2576
rect 13537 2544 16871 2546
rect 13537 2488 13542 2544
rect 13598 2488 16871 2544
rect 13537 2486 16871 2488
rect 13537 2483 13603 2486
rect 16071 2456 16871 2486
rect 5820 2208 6140 2209
rect 5820 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6140 2208
rect 5820 2143 6140 2144
rect 10696 2208 11016 2209
rect 10696 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11016 2208
rect 10696 2143 11016 2144
<< via3 >>
rect 5828 16348 5892 16352
rect 5828 16292 5832 16348
rect 5832 16292 5888 16348
rect 5888 16292 5892 16348
rect 5828 16288 5892 16292
rect 5908 16348 5972 16352
rect 5908 16292 5912 16348
rect 5912 16292 5968 16348
rect 5968 16292 5972 16348
rect 5908 16288 5972 16292
rect 5988 16348 6052 16352
rect 5988 16292 5992 16348
rect 5992 16292 6048 16348
rect 6048 16292 6052 16348
rect 5988 16288 6052 16292
rect 6068 16348 6132 16352
rect 6068 16292 6072 16348
rect 6072 16292 6128 16348
rect 6128 16292 6132 16348
rect 6068 16288 6132 16292
rect 10704 16348 10768 16352
rect 10704 16292 10708 16348
rect 10708 16292 10764 16348
rect 10764 16292 10768 16348
rect 10704 16288 10768 16292
rect 10784 16348 10848 16352
rect 10784 16292 10788 16348
rect 10788 16292 10844 16348
rect 10844 16292 10848 16348
rect 10784 16288 10848 16292
rect 10864 16348 10928 16352
rect 10864 16292 10868 16348
rect 10868 16292 10924 16348
rect 10924 16292 10928 16348
rect 10864 16288 10928 16292
rect 10944 16348 11008 16352
rect 10944 16292 10948 16348
rect 10948 16292 11004 16348
rect 11004 16292 11008 16348
rect 10944 16288 11008 16292
rect 3390 15804 3454 15808
rect 3390 15748 3394 15804
rect 3394 15748 3450 15804
rect 3450 15748 3454 15804
rect 3390 15744 3454 15748
rect 3470 15804 3534 15808
rect 3470 15748 3474 15804
rect 3474 15748 3530 15804
rect 3530 15748 3534 15804
rect 3470 15744 3534 15748
rect 3550 15804 3614 15808
rect 3550 15748 3554 15804
rect 3554 15748 3610 15804
rect 3610 15748 3614 15804
rect 3550 15744 3614 15748
rect 3630 15804 3694 15808
rect 3630 15748 3634 15804
rect 3634 15748 3690 15804
rect 3690 15748 3694 15804
rect 3630 15744 3694 15748
rect 8266 15804 8330 15808
rect 8266 15748 8270 15804
rect 8270 15748 8326 15804
rect 8326 15748 8330 15804
rect 8266 15744 8330 15748
rect 8346 15804 8410 15808
rect 8346 15748 8350 15804
rect 8350 15748 8406 15804
rect 8406 15748 8410 15804
rect 8346 15744 8410 15748
rect 8426 15804 8490 15808
rect 8426 15748 8430 15804
rect 8430 15748 8486 15804
rect 8486 15748 8490 15804
rect 8426 15744 8490 15748
rect 8506 15804 8570 15808
rect 8506 15748 8510 15804
rect 8510 15748 8566 15804
rect 8566 15748 8570 15804
rect 8506 15744 8570 15748
rect 13142 15804 13206 15808
rect 13142 15748 13146 15804
rect 13146 15748 13202 15804
rect 13202 15748 13206 15804
rect 13142 15744 13206 15748
rect 13222 15804 13286 15808
rect 13222 15748 13226 15804
rect 13226 15748 13282 15804
rect 13282 15748 13286 15804
rect 13222 15744 13286 15748
rect 13302 15804 13366 15808
rect 13302 15748 13306 15804
rect 13306 15748 13362 15804
rect 13362 15748 13366 15804
rect 13302 15744 13366 15748
rect 13382 15804 13446 15808
rect 13382 15748 13386 15804
rect 13386 15748 13442 15804
rect 13442 15748 13446 15804
rect 13382 15744 13446 15748
rect 5828 15260 5892 15264
rect 5828 15204 5832 15260
rect 5832 15204 5888 15260
rect 5888 15204 5892 15260
rect 5828 15200 5892 15204
rect 5908 15260 5972 15264
rect 5908 15204 5912 15260
rect 5912 15204 5968 15260
rect 5968 15204 5972 15260
rect 5908 15200 5972 15204
rect 5988 15260 6052 15264
rect 5988 15204 5992 15260
rect 5992 15204 6048 15260
rect 6048 15204 6052 15260
rect 5988 15200 6052 15204
rect 6068 15260 6132 15264
rect 6068 15204 6072 15260
rect 6072 15204 6128 15260
rect 6128 15204 6132 15260
rect 6068 15200 6132 15204
rect 10704 15260 10768 15264
rect 10704 15204 10708 15260
rect 10708 15204 10764 15260
rect 10764 15204 10768 15260
rect 10704 15200 10768 15204
rect 10784 15260 10848 15264
rect 10784 15204 10788 15260
rect 10788 15204 10844 15260
rect 10844 15204 10848 15260
rect 10784 15200 10848 15204
rect 10864 15260 10928 15264
rect 10864 15204 10868 15260
rect 10868 15204 10924 15260
rect 10924 15204 10928 15260
rect 10864 15200 10928 15204
rect 10944 15260 11008 15264
rect 10944 15204 10948 15260
rect 10948 15204 11004 15260
rect 11004 15204 11008 15260
rect 10944 15200 11008 15204
rect 3390 14716 3454 14720
rect 3390 14660 3394 14716
rect 3394 14660 3450 14716
rect 3450 14660 3454 14716
rect 3390 14656 3454 14660
rect 3470 14716 3534 14720
rect 3470 14660 3474 14716
rect 3474 14660 3530 14716
rect 3530 14660 3534 14716
rect 3470 14656 3534 14660
rect 3550 14716 3614 14720
rect 3550 14660 3554 14716
rect 3554 14660 3610 14716
rect 3610 14660 3614 14716
rect 3550 14656 3614 14660
rect 3630 14716 3694 14720
rect 3630 14660 3634 14716
rect 3634 14660 3690 14716
rect 3690 14660 3694 14716
rect 3630 14656 3694 14660
rect 8266 14716 8330 14720
rect 8266 14660 8270 14716
rect 8270 14660 8326 14716
rect 8326 14660 8330 14716
rect 8266 14656 8330 14660
rect 8346 14716 8410 14720
rect 8346 14660 8350 14716
rect 8350 14660 8406 14716
rect 8406 14660 8410 14716
rect 8346 14656 8410 14660
rect 8426 14716 8490 14720
rect 8426 14660 8430 14716
rect 8430 14660 8486 14716
rect 8486 14660 8490 14716
rect 8426 14656 8490 14660
rect 8506 14716 8570 14720
rect 8506 14660 8510 14716
rect 8510 14660 8566 14716
rect 8566 14660 8570 14716
rect 8506 14656 8570 14660
rect 13142 14716 13206 14720
rect 13142 14660 13146 14716
rect 13146 14660 13202 14716
rect 13202 14660 13206 14716
rect 13142 14656 13206 14660
rect 13222 14716 13286 14720
rect 13222 14660 13226 14716
rect 13226 14660 13282 14716
rect 13282 14660 13286 14716
rect 13222 14656 13286 14660
rect 13302 14716 13366 14720
rect 13302 14660 13306 14716
rect 13306 14660 13362 14716
rect 13362 14660 13366 14716
rect 13302 14656 13366 14660
rect 13382 14716 13446 14720
rect 13382 14660 13386 14716
rect 13386 14660 13442 14716
rect 13442 14660 13446 14716
rect 13382 14656 13446 14660
rect 5828 14172 5892 14176
rect 5828 14116 5832 14172
rect 5832 14116 5888 14172
rect 5888 14116 5892 14172
rect 5828 14112 5892 14116
rect 5908 14172 5972 14176
rect 5908 14116 5912 14172
rect 5912 14116 5968 14172
rect 5968 14116 5972 14172
rect 5908 14112 5972 14116
rect 5988 14172 6052 14176
rect 5988 14116 5992 14172
rect 5992 14116 6048 14172
rect 6048 14116 6052 14172
rect 5988 14112 6052 14116
rect 6068 14172 6132 14176
rect 6068 14116 6072 14172
rect 6072 14116 6128 14172
rect 6128 14116 6132 14172
rect 6068 14112 6132 14116
rect 10704 14172 10768 14176
rect 10704 14116 10708 14172
rect 10708 14116 10764 14172
rect 10764 14116 10768 14172
rect 10704 14112 10768 14116
rect 10784 14172 10848 14176
rect 10784 14116 10788 14172
rect 10788 14116 10844 14172
rect 10844 14116 10848 14172
rect 10784 14112 10848 14116
rect 10864 14172 10928 14176
rect 10864 14116 10868 14172
rect 10868 14116 10924 14172
rect 10924 14116 10928 14172
rect 10864 14112 10928 14116
rect 10944 14172 11008 14176
rect 10944 14116 10948 14172
rect 10948 14116 11004 14172
rect 11004 14116 11008 14172
rect 10944 14112 11008 14116
rect 3390 13628 3454 13632
rect 3390 13572 3394 13628
rect 3394 13572 3450 13628
rect 3450 13572 3454 13628
rect 3390 13568 3454 13572
rect 3470 13628 3534 13632
rect 3470 13572 3474 13628
rect 3474 13572 3530 13628
rect 3530 13572 3534 13628
rect 3470 13568 3534 13572
rect 3550 13628 3614 13632
rect 3550 13572 3554 13628
rect 3554 13572 3610 13628
rect 3610 13572 3614 13628
rect 3550 13568 3614 13572
rect 3630 13628 3694 13632
rect 3630 13572 3634 13628
rect 3634 13572 3690 13628
rect 3690 13572 3694 13628
rect 3630 13568 3694 13572
rect 8266 13628 8330 13632
rect 8266 13572 8270 13628
rect 8270 13572 8326 13628
rect 8326 13572 8330 13628
rect 8266 13568 8330 13572
rect 8346 13628 8410 13632
rect 8346 13572 8350 13628
rect 8350 13572 8406 13628
rect 8406 13572 8410 13628
rect 8346 13568 8410 13572
rect 8426 13628 8490 13632
rect 8426 13572 8430 13628
rect 8430 13572 8486 13628
rect 8486 13572 8490 13628
rect 8426 13568 8490 13572
rect 8506 13628 8570 13632
rect 8506 13572 8510 13628
rect 8510 13572 8566 13628
rect 8566 13572 8570 13628
rect 8506 13568 8570 13572
rect 13142 13628 13206 13632
rect 13142 13572 13146 13628
rect 13146 13572 13202 13628
rect 13202 13572 13206 13628
rect 13142 13568 13206 13572
rect 13222 13628 13286 13632
rect 13222 13572 13226 13628
rect 13226 13572 13282 13628
rect 13282 13572 13286 13628
rect 13222 13568 13286 13572
rect 13302 13628 13366 13632
rect 13302 13572 13306 13628
rect 13306 13572 13362 13628
rect 13362 13572 13366 13628
rect 13302 13568 13366 13572
rect 13382 13628 13446 13632
rect 13382 13572 13386 13628
rect 13386 13572 13442 13628
rect 13442 13572 13446 13628
rect 13382 13568 13446 13572
rect 5828 13084 5892 13088
rect 5828 13028 5832 13084
rect 5832 13028 5888 13084
rect 5888 13028 5892 13084
rect 5828 13024 5892 13028
rect 5908 13084 5972 13088
rect 5908 13028 5912 13084
rect 5912 13028 5968 13084
rect 5968 13028 5972 13084
rect 5908 13024 5972 13028
rect 5988 13084 6052 13088
rect 5988 13028 5992 13084
rect 5992 13028 6048 13084
rect 6048 13028 6052 13084
rect 5988 13024 6052 13028
rect 6068 13084 6132 13088
rect 6068 13028 6072 13084
rect 6072 13028 6128 13084
rect 6128 13028 6132 13084
rect 6068 13024 6132 13028
rect 10704 13084 10768 13088
rect 10704 13028 10708 13084
rect 10708 13028 10764 13084
rect 10764 13028 10768 13084
rect 10704 13024 10768 13028
rect 10784 13084 10848 13088
rect 10784 13028 10788 13084
rect 10788 13028 10844 13084
rect 10844 13028 10848 13084
rect 10784 13024 10848 13028
rect 10864 13084 10928 13088
rect 10864 13028 10868 13084
rect 10868 13028 10924 13084
rect 10924 13028 10928 13084
rect 10864 13024 10928 13028
rect 10944 13084 11008 13088
rect 10944 13028 10948 13084
rect 10948 13028 11004 13084
rect 11004 13028 11008 13084
rect 10944 13024 11008 13028
rect 3390 12540 3454 12544
rect 3390 12484 3394 12540
rect 3394 12484 3450 12540
rect 3450 12484 3454 12540
rect 3390 12480 3454 12484
rect 3470 12540 3534 12544
rect 3470 12484 3474 12540
rect 3474 12484 3530 12540
rect 3530 12484 3534 12540
rect 3470 12480 3534 12484
rect 3550 12540 3614 12544
rect 3550 12484 3554 12540
rect 3554 12484 3610 12540
rect 3610 12484 3614 12540
rect 3550 12480 3614 12484
rect 3630 12540 3694 12544
rect 3630 12484 3634 12540
rect 3634 12484 3690 12540
rect 3690 12484 3694 12540
rect 3630 12480 3694 12484
rect 8266 12540 8330 12544
rect 8266 12484 8270 12540
rect 8270 12484 8326 12540
rect 8326 12484 8330 12540
rect 8266 12480 8330 12484
rect 8346 12540 8410 12544
rect 8346 12484 8350 12540
rect 8350 12484 8406 12540
rect 8406 12484 8410 12540
rect 8346 12480 8410 12484
rect 8426 12540 8490 12544
rect 8426 12484 8430 12540
rect 8430 12484 8486 12540
rect 8486 12484 8490 12540
rect 8426 12480 8490 12484
rect 8506 12540 8570 12544
rect 8506 12484 8510 12540
rect 8510 12484 8566 12540
rect 8566 12484 8570 12540
rect 8506 12480 8570 12484
rect 13142 12540 13206 12544
rect 13142 12484 13146 12540
rect 13146 12484 13202 12540
rect 13202 12484 13206 12540
rect 13142 12480 13206 12484
rect 13222 12540 13286 12544
rect 13222 12484 13226 12540
rect 13226 12484 13282 12540
rect 13282 12484 13286 12540
rect 13222 12480 13286 12484
rect 13302 12540 13366 12544
rect 13302 12484 13306 12540
rect 13306 12484 13362 12540
rect 13362 12484 13366 12540
rect 13302 12480 13366 12484
rect 13382 12540 13446 12544
rect 13382 12484 13386 12540
rect 13386 12484 13442 12540
rect 13442 12484 13446 12540
rect 13382 12480 13446 12484
rect 5828 11996 5892 12000
rect 5828 11940 5832 11996
rect 5832 11940 5888 11996
rect 5888 11940 5892 11996
rect 5828 11936 5892 11940
rect 5908 11996 5972 12000
rect 5908 11940 5912 11996
rect 5912 11940 5968 11996
rect 5968 11940 5972 11996
rect 5908 11936 5972 11940
rect 5988 11996 6052 12000
rect 5988 11940 5992 11996
rect 5992 11940 6048 11996
rect 6048 11940 6052 11996
rect 5988 11936 6052 11940
rect 6068 11996 6132 12000
rect 6068 11940 6072 11996
rect 6072 11940 6128 11996
rect 6128 11940 6132 11996
rect 6068 11936 6132 11940
rect 10704 11996 10768 12000
rect 10704 11940 10708 11996
rect 10708 11940 10764 11996
rect 10764 11940 10768 11996
rect 10704 11936 10768 11940
rect 10784 11996 10848 12000
rect 10784 11940 10788 11996
rect 10788 11940 10844 11996
rect 10844 11940 10848 11996
rect 10784 11936 10848 11940
rect 10864 11996 10928 12000
rect 10864 11940 10868 11996
rect 10868 11940 10924 11996
rect 10924 11940 10928 11996
rect 10864 11936 10928 11940
rect 10944 11996 11008 12000
rect 10944 11940 10948 11996
rect 10948 11940 11004 11996
rect 11004 11940 11008 11996
rect 10944 11936 11008 11940
rect 3390 11452 3454 11456
rect 3390 11396 3394 11452
rect 3394 11396 3450 11452
rect 3450 11396 3454 11452
rect 3390 11392 3454 11396
rect 3470 11452 3534 11456
rect 3470 11396 3474 11452
rect 3474 11396 3530 11452
rect 3530 11396 3534 11452
rect 3470 11392 3534 11396
rect 3550 11452 3614 11456
rect 3550 11396 3554 11452
rect 3554 11396 3610 11452
rect 3610 11396 3614 11452
rect 3550 11392 3614 11396
rect 3630 11452 3694 11456
rect 3630 11396 3634 11452
rect 3634 11396 3690 11452
rect 3690 11396 3694 11452
rect 3630 11392 3694 11396
rect 8266 11452 8330 11456
rect 8266 11396 8270 11452
rect 8270 11396 8326 11452
rect 8326 11396 8330 11452
rect 8266 11392 8330 11396
rect 8346 11452 8410 11456
rect 8346 11396 8350 11452
rect 8350 11396 8406 11452
rect 8406 11396 8410 11452
rect 8346 11392 8410 11396
rect 8426 11452 8490 11456
rect 8426 11396 8430 11452
rect 8430 11396 8486 11452
rect 8486 11396 8490 11452
rect 8426 11392 8490 11396
rect 8506 11452 8570 11456
rect 8506 11396 8510 11452
rect 8510 11396 8566 11452
rect 8566 11396 8570 11452
rect 8506 11392 8570 11396
rect 13142 11452 13206 11456
rect 13142 11396 13146 11452
rect 13146 11396 13202 11452
rect 13202 11396 13206 11452
rect 13142 11392 13206 11396
rect 13222 11452 13286 11456
rect 13222 11396 13226 11452
rect 13226 11396 13282 11452
rect 13282 11396 13286 11452
rect 13222 11392 13286 11396
rect 13302 11452 13366 11456
rect 13302 11396 13306 11452
rect 13306 11396 13362 11452
rect 13362 11396 13366 11452
rect 13302 11392 13366 11396
rect 13382 11452 13446 11456
rect 13382 11396 13386 11452
rect 13386 11396 13442 11452
rect 13442 11396 13446 11452
rect 13382 11392 13446 11396
rect 5828 10908 5892 10912
rect 5828 10852 5832 10908
rect 5832 10852 5888 10908
rect 5888 10852 5892 10908
rect 5828 10848 5892 10852
rect 5908 10908 5972 10912
rect 5908 10852 5912 10908
rect 5912 10852 5968 10908
rect 5968 10852 5972 10908
rect 5908 10848 5972 10852
rect 5988 10908 6052 10912
rect 5988 10852 5992 10908
rect 5992 10852 6048 10908
rect 6048 10852 6052 10908
rect 5988 10848 6052 10852
rect 6068 10908 6132 10912
rect 6068 10852 6072 10908
rect 6072 10852 6128 10908
rect 6128 10852 6132 10908
rect 6068 10848 6132 10852
rect 10704 10908 10768 10912
rect 10704 10852 10708 10908
rect 10708 10852 10764 10908
rect 10764 10852 10768 10908
rect 10704 10848 10768 10852
rect 10784 10908 10848 10912
rect 10784 10852 10788 10908
rect 10788 10852 10844 10908
rect 10844 10852 10848 10908
rect 10784 10848 10848 10852
rect 10864 10908 10928 10912
rect 10864 10852 10868 10908
rect 10868 10852 10924 10908
rect 10924 10852 10928 10908
rect 10864 10848 10928 10852
rect 10944 10908 11008 10912
rect 10944 10852 10948 10908
rect 10948 10852 11004 10908
rect 11004 10852 11008 10908
rect 10944 10848 11008 10852
rect 3390 10364 3454 10368
rect 3390 10308 3394 10364
rect 3394 10308 3450 10364
rect 3450 10308 3454 10364
rect 3390 10304 3454 10308
rect 3470 10364 3534 10368
rect 3470 10308 3474 10364
rect 3474 10308 3530 10364
rect 3530 10308 3534 10364
rect 3470 10304 3534 10308
rect 3550 10364 3614 10368
rect 3550 10308 3554 10364
rect 3554 10308 3610 10364
rect 3610 10308 3614 10364
rect 3550 10304 3614 10308
rect 3630 10364 3694 10368
rect 3630 10308 3634 10364
rect 3634 10308 3690 10364
rect 3690 10308 3694 10364
rect 3630 10304 3694 10308
rect 8266 10364 8330 10368
rect 8266 10308 8270 10364
rect 8270 10308 8326 10364
rect 8326 10308 8330 10364
rect 8266 10304 8330 10308
rect 8346 10364 8410 10368
rect 8346 10308 8350 10364
rect 8350 10308 8406 10364
rect 8406 10308 8410 10364
rect 8346 10304 8410 10308
rect 8426 10364 8490 10368
rect 8426 10308 8430 10364
rect 8430 10308 8486 10364
rect 8486 10308 8490 10364
rect 8426 10304 8490 10308
rect 8506 10364 8570 10368
rect 8506 10308 8510 10364
rect 8510 10308 8566 10364
rect 8566 10308 8570 10364
rect 8506 10304 8570 10308
rect 13142 10364 13206 10368
rect 13142 10308 13146 10364
rect 13146 10308 13202 10364
rect 13202 10308 13206 10364
rect 13142 10304 13206 10308
rect 13222 10364 13286 10368
rect 13222 10308 13226 10364
rect 13226 10308 13282 10364
rect 13282 10308 13286 10364
rect 13222 10304 13286 10308
rect 13302 10364 13366 10368
rect 13302 10308 13306 10364
rect 13306 10308 13362 10364
rect 13362 10308 13366 10364
rect 13302 10304 13366 10308
rect 13382 10364 13446 10368
rect 13382 10308 13386 10364
rect 13386 10308 13442 10364
rect 13442 10308 13446 10364
rect 13382 10304 13446 10308
rect 5828 9820 5892 9824
rect 5828 9764 5832 9820
rect 5832 9764 5888 9820
rect 5888 9764 5892 9820
rect 5828 9760 5892 9764
rect 5908 9820 5972 9824
rect 5908 9764 5912 9820
rect 5912 9764 5968 9820
rect 5968 9764 5972 9820
rect 5908 9760 5972 9764
rect 5988 9820 6052 9824
rect 5988 9764 5992 9820
rect 5992 9764 6048 9820
rect 6048 9764 6052 9820
rect 5988 9760 6052 9764
rect 6068 9820 6132 9824
rect 6068 9764 6072 9820
rect 6072 9764 6128 9820
rect 6128 9764 6132 9820
rect 6068 9760 6132 9764
rect 10704 9820 10768 9824
rect 10704 9764 10708 9820
rect 10708 9764 10764 9820
rect 10764 9764 10768 9820
rect 10704 9760 10768 9764
rect 10784 9820 10848 9824
rect 10784 9764 10788 9820
rect 10788 9764 10844 9820
rect 10844 9764 10848 9820
rect 10784 9760 10848 9764
rect 10864 9820 10928 9824
rect 10864 9764 10868 9820
rect 10868 9764 10924 9820
rect 10924 9764 10928 9820
rect 10864 9760 10928 9764
rect 10944 9820 11008 9824
rect 10944 9764 10948 9820
rect 10948 9764 11004 9820
rect 11004 9764 11008 9820
rect 10944 9760 11008 9764
rect 3390 9276 3454 9280
rect 3390 9220 3394 9276
rect 3394 9220 3450 9276
rect 3450 9220 3454 9276
rect 3390 9216 3454 9220
rect 3470 9276 3534 9280
rect 3470 9220 3474 9276
rect 3474 9220 3530 9276
rect 3530 9220 3534 9276
rect 3470 9216 3534 9220
rect 3550 9276 3614 9280
rect 3550 9220 3554 9276
rect 3554 9220 3610 9276
rect 3610 9220 3614 9276
rect 3550 9216 3614 9220
rect 3630 9276 3694 9280
rect 3630 9220 3634 9276
rect 3634 9220 3690 9276
rect 3690 9220 3694 9276
rect 3630 9216 3694 9220
rect 8266 9276 8330 9280
rect 8266 9220 8270 9276
rect 8270 9220 8326 9276
rect 8326 9220 8330 9276
rect 8266 9216 8330 9220
rect 8346 9276 8410 9280
rect 8346 9220 8350 9276
rect 8350 9220 8406 9276
rect 8406 9220 8410 9276
rect 8346 9216 8410 9220
rect 8426 9276 8490 9280
rect 8426 9220 8430 9276
rect 8430 9220 8486 9276
rect 8486 9220 8490 9276
rect 8426 9216 8490 9220
rect 8506 9276 8570 9280
rect 8506 9220 8510 9276
rect 8510 9220 8566 9276
rect 8566 9220 8570 9276
rect 8506 9216 8570 9220
rect 13142 9276 13206 9280
rect 13142 9220 13146 9276
rect 13146 9220 13202 9276
rect 13202 9220 13206 9276
rect 13142 9216 13206 9220
rect 13222 9276 13286 9280
rect 13222 9220 13226 9276
rect 13226 9220 13282 9276
rect 13282 9220 13286 9276
rect 13222 9216 13286 9220
rect 13302 9276 13366 9280
rect 13302 9220 13306 9276
rect 13306 9220 13362 9276
rect 13362 9220 13366 9276
rect 13302 9216 13366 9220
rect 13382 9276 13446 9280
rect 13382 9220 13386 9276
rect 13386 9220 13442 9276
rect 13442 9220 13446 9276
rect 13382 9216 13446 9220
rect 5828 8732 5892 8736
rect 5828 8676 5832 8732
rect 5832 8676 5888 8732
rect 5888 8676 5892 8732
rect 5828 8672 5892 8676
rect 5908 8732 5972 8736
rect 5908 8676 5912 8732
rect 5912 8676 5968 8732
rect 5968 8676 5972 8732
rect 5908 8672 5972 8676
rect 5988 8732 6052 8736
rect 5988 8676 5992 8732
rect 5992 8676 6048 8732
rect 6048 8676 6052 8732
rect 5988 8672 6052 8676
rect 6068 8732 6132 8736
rect 6068 8676 6072 8732
rect 6072 8676 6128 8732
rect 6128 8676 6132 8732
rect 6068 8672 6132 8676
rect 10704 8732 10768 8736
rect 10704 8676 10708 8732
rect 10708 8676 10764 8732
rect 10764 8676 10768 8732
rect 10704 8672 10768 8676
rect 10784 8732 10848 8736
rect 10784 8676 10788 8732
rect 10788 8676 10844 8732
rect 10844 8676 10848 8732
rect 10784 8672 10848 8676
rect 10864 8732 10928 8736
rect 10864 8676 10868 8732
rect 10868 8676 10924 8732
rect 10924 8676 10928 8732
rect 10864 8672 10928 8676
rect 10944 8732 11008 8736
rect 10944 8676 10948 8732
rect 10948 8676 11004 8732
rect 11004 8676 11008 8732
rect 10944 8672 11008 8676
rect 3390 8188 3454 8192
rect 3390 8132 3394 8188
rect 3394 8132 3450 8188
rect 3450 8132 3454 8188
rect 3390 8128 3454 8132
rect 3470 8188 3534 8192
rect 3470 8132 3474 8188
rect 3474 8132 3530 8188
rect 3530 8132 3534 8188
rect 3470 8128 3534 8132
rect 3550 8188 3614 8192
rect 3550 8132 3554 8188
rect 3554 8132 3610 8188
rect 3610 8132 3614 8188
rect 3550 8128 3614 8132
rect 3630 8188 3694 8192
rect 3630 8132 3634 8188
rect 3634 8132 3690 8188
rect 3690 8132 3694 8188
rect 3630 8128 3694 8132
rect 8266 8188 8330 8192
rect 8266 8132 8270 8188
rect 8270 8132 8326 8188
rect 8326 8132 8330 8188
rect 8266 8128 8330 8132
rect 8346 8188 8410 8192
rect 8346 8132 8350 8188
rect 8350 8132 8406 8188
rect 8406 8132 8410 8188
rect 8346 8128 8410 8132
rect 8426 8188 8490 8192
rect 8426 8132 8430 8188
rect 8430 8132 8486 8188
rect 8486 8132 8490 8188
rect 8426 8128 8490 8132
rect 8506 8188 8570 8192
rect 8506 8132 8510 8188
rect 8510 8132 8566 8188
rect 8566 8132 8570 8188
rect 8506 8128 8570 8132
rect 13142 8188 13206 8192
rect 13142 8132 13146 8188
rect 13146 8132 13202 8188
rect 13202 8132 13206 8188
rect 13142 8128 13206 8132
rect 13222 8188 13286 8192
rect 13222 8132 13226 8188
rect 13226 8132 13282 8188
rect 13282 8132 13286 8188
rect 13222 8128 13286 8132
rect 13302 8188 13366 8192
rect 13302 8132 13306 8188
rect 13306 8132 13362 8188
rect 13362 8132 13366 8188
rect 13302 8128 13366 8132
rect 13382 8188 13446 8192
rect 13382 8132 13386 8188
rect 13386 8132 13442 8188
rect 13442 8132 13446 8188
rect 13382 8128 13446 8132
rect 5828 7644 5892 7648
rect 5828 7588 5832 7644
rect 5832 7588 5888 7644
rect 5888 7588 5892 7644
rect 5828 7584 5892 7588
rect 5908 7644 5972 7648
rect 5908 7588 5912 7644
rect 5912 7588 5968 7644
rect 5968 7588 5972 7644
rect 5908 7584 5972 7588
rect 5988 7644 6052 7648
rect 5988 7588 5992 7644
rect 5992 7588 6048 7644
rect 6048 7588 6052 7644
rect 5988 7584 6052 7588
rect 6068 7644 6132 7648
rect 6068 7588 6072 7644
rect 6072 7588 6128 7644
rect 6128 7588 6132 7644
rect 6068 7584 6132 7588
rect 10704 7644 10768 7648
rect 10704 7588 10708 7644
rect 10708 7588 10764 7644
rect 10764 7588 10768 7644
rect 10704 7584 10768 7588
rect 10784 7644 10848 7648
rect 10784 7588 10788 7644
rect 10788 7588 10844 7644
rect 10844 7588 10848 7644
rect 10784 7584 10848 7588
rect 10864 7644 10928 7648
rect 10864 7588 10868 7644
rect 10868 7588 10924 7644
rect 10924 7588 10928 7644
rect 10864 7584 10928 7588
rect 10944 7644 11008 7648
rect 10944 7588 10948 7644
rect 10948 7588 11004 7644
rect 11004 7588 11008 7644
rect 10944 7584 11008 7588
rect 3390 7100 3454 7104
rect 3390 7044 3394 7100
rect 3394 7044 3450 7100
rect 3450 7044 3454 7100
rect 3390 7040 3454 7044
rect 3470 7100 3534 7104
rect 3470 7044 3474 7100
rect 3474 7044 3530 7100
rect 3530 7044 3534 7100
rect 3470 7040 3534 7044
rect 3550 7100 3614 7104
rect 3550 7044 3554 7100
rect 3554 7044 3610 7100
rect 3610 7044 3614 7100
rect 3550 7040 3614 7044
rect 3630 7100 3694 7104
rect 3630 7044 3634 7100
rect 3634 7044 3690 7100
rect 3690 7044 3694 7100
rect 3630 7040 3694 7044
rect 8266 7100 8330 7104
rect 8266 7044 8270 7100
rect 8270 7044 8326 7100
rect 8326 7044 8330 7100
rect 8266 7040 8330 7044
rect 8346 7100 8410 7104
rect 8346 7044 8350 7100
rect 8350 7044 8406 7100
rect 8406 7044 8410 7100
rect 8346 7040 8410 7044
rect 8426 7100 8490 7104
rect 8426 7044 8430 7100
rect 8430 7044 8486 7100
rect 8486 7044 8490 7100
rect 8426 7040 8490 7044
rect 8506 7100 8570 7104
rect 8506 7044 8510 7100
rect 8510 7044 8566 7100
rect 8566 7044 8570 7100
rect 8506 7040 8570 7044
rect 13142 7100 13206 7104
rect 13142 7044 13146 7100
rect 13146 7044 13202 7100
rect 13202 7044 13206 7100
rect 13142 7040 13206 7044
rect 13222 7100 13286 7104
rect 13222 7044 13226 7100
rect 13226 7044 13282 7100
rect 13282 7044 13286 7100
rect 13222 7040 13286 7044
rect 13302 7100 13366 7104
rect 13302 7044 13306 7100
rect 13306 7044 13362 7100
rect 13362 7044 13366 7100
rect 13302 7040 13366 7044
rect 13382 7100 13446 7104
rect 13382 7044 13386 7100
rect 13386 7044 13442 7100
rect 13442 7044 13446 7100
rect 13382 7040 13446 7044
rect 5828 6556 5892 6560
rect 5828 6500 5832 6556
rect 5832 6500 5888 6556
rect 5888 6500 5892 6556
rect 5828 6496 5892 6500
rect 5908 6556 5972 6560
rect 5908 6500 5912 6556
rect 5912 6500 5968 6556
rect 5968 6500 5972 6556
rect 5908 6496 5972 6500
rect 5988 6556 6052 6560
rect 5988 6500 5992 6556
rect 5992 6500 6048 6556
rect 6048 6500 6052 6556
rect 5988 6496 6052 6500
rect 6068 6556 6132 6560
rect 6068 6500 6072 6556
rect 6072 6500 6128 6556
rect 6128 6500 6132 6556
rect 6068 6496 6132 6500
rect 10704 6556 10768 6560
rect 10704 6500 10708 6556
rect 10708 6500 10764 6556
rect 10764 6500 10768 6556
rect 10704 6496 10768 6500
rect 10784 6556 10848 6560
rect 10784 6500 10788 6556
rect 10788 6500 10844 6556
rect 10844 6500 10848 6556
rect 10784 6496 10848 6500
rect 10864 6556 10928 6560
rect 10864 6500 10868 6556
rect 10868 6500 10924 6556
rect 10924 6500 10928 6556
rect 10864 6496 10928 6500
rect 10944 6556 11008 6560
rect 10944 6500 10948 6556
rect 10948 6500 11004 6556
rect 11004 6500 11008 6556
rect 10944 6496 11008 6500
rect 3390 6012 3454 6016
rect 3390 5956 3394 6012
rect 3394 5956 3450 6012
rect 3450 5956 3454 6012
rect 3390 5952 3454 5956
rect 3470 6012 3534 6016
rect 3470 5956 3474 6012
rect 3474 5956 3530 6012
rect 3530 5956 3534 6012
rect 3470 5952 3534 5956
rect 3550 6012 3614 6016
rect 3550 5956 3554 6012
rect 3554 5956 3610 6012
rect 3610 5956 3614 6012
rect 3550 5952 3614 5956
rect 3630 6012 3694 6016
rect 3630 5956 3634 6012
rect 3634 5956 3690 6012
rect 3690 5956 3694 6012
rect 3630 5952 3694 5956
rect 8266 6012 8330 6016
rect 8266 5956 8270 6012
rect 8270 5956 8326 6012
rect 8326 5956 8330 6012
rect 8266 5952 8330 5956
rect 8346 6012 8410 6016
rect 8346 5956 8350 6012
rect 8350 5956 8406 6012
rect 8406 5956 8410 6012
rect 8346 5952 8410 5956
rect 8426 6012 8490 6016
rect 8426 5956 8430 6012
rect 8430 5956 8486 6012
rect 8486 5956 8490 6012
rect 8426 5952 8490 5956
rect 8506 6012 8570 6016
rect 8506 5956 8510 6012
rect 8510 5956 8566 6012
rect 8566 5956 8570 6012
rect 8506 5952 8570 5956
rect 13142 6012 13206 6016
rect 13142 5956 13146 6012
rect 13146 5956 13202 6012
rect 13202 5956 13206 6012
rect 13142 5952 13206 5956
rect 13222 6012 13286 6016
rect 13222 5956 13226 6012
rect 13226 5956 13282 6012
rect 13282 5956 13286 6012
rect 13222 5952 13286 5956
rect 13302 6012 13366 6016
rect 13302 5956 13306 6012
rect 13306 5956 13362 6012
rect 13362 5956 13366 6012
rect 13302 5952 13366 5956
rect 13382 6012 13446 6016
rect 13382 5956 13386 6012
rect 13386 5956 13442 6012
rect 13442 5956 13446 6012
rect 13382 5952 13446 5956
rect 5828 5468 5892 5472
rect 5828 5412 5832 5468
rect 5832 5412 5888 5468
rect 5888 5412 5892 5468
rect 5828 5408 5892 5412
rect 5908 5468 5972 5472
rect 5908 5412 5912 5468
rect 5912 5412 5968 5468
rect 5968 5412 5972 5468
rect 5908 5408 5972 5412
rect 5988 5468 6052 5472
rect 5988 5412 5992 5468
rect 5992 5412 6048 5468
rect 6048 5412 6052 5468
rect 5988 5408 6052 5412
rect 6068 5468 6132 5472
rect 6068 5412 6072 5468
rect 6072 5412 6128 5468
rect 6128 5412 6132 5468
rect 6068 5408 6132 5412
rect 10704 5468 10768 5472
rect 10704 5412 10708 5468
rect 10708 5412 10764 5468
rect 10764 5412 10768 5468
rect 10704 5408 10768 5412
rect 10784 5468 10848 5472
rect 10784 5412 10788 5468
rect 10788 5412 10844 5468
rect 10844 5412 10848 5468
rect 10784 5408 10848 5412
rect 10864 5468 10928 5472
rect 10864 5412 10868 5468
rect 10868 5412 10924 5468
rect 10924 5412 10928 5468
rect 10864 5408 10928 5412
rect 10944 5468 11008 5472
rect 10944 5412 10948 5468
rect 10948 5412 11004 5468
rect 11004 5412 11008 5468
rect 10944 5408 11008 5412
rect 3390 4924 3454 4928
rect 3390 4868 3394 4924
rect 3394 4868 3450 4924
rect 3450 4868 3454 4924
rect 3390 4864 3454 4868
rect 3470 4924 3534 4928
rect 3470 4868 3474 4924
rect 3474 4868 3530 4924
rect 3530 4868 3534 4924
rect 3470 4864 3534 4868
rect 3550 4924 3614 4928
rect 3550 4868 3554 4924
rect 3554 4868 3610 4924
rect 3610 4868 3614 4924
rect 3550 4864 3614 4868
rect 3630 4924 3694 4928
rect 3630 4868 3634 4924
rect 3634 4868 3690 4924
rect 3690 4868 3694 4924
rect 3630 4864 3694 4868
rect 8266 4924 8330 4928
rect 8266 4868 8270 4924
rect 8270 4868 8326 4924
rect 8326 4868 8330 4924
rect 8266 4864 8330 4868
rect 8346 4924 8410 4928
rect 8346 4868 8350 4924
rect 8350 4868 8406 4924
rect 8406 4868 8410 4924
rect 8346 4864 8410 4868
rect 8426 4924 8490 4928
rect 8426 4868 8430 4924
rect 8430 4868 8486 4924
rect 8486 4868 8490 4924
rect 8426 4864 8490 4868
rect 8506 4924 8570 4928
rect 8506 4868 8510 4924
rect 8510 4868 8566 4924
rect 8566 4868 8570 4924
rect 8506 4864 8570 4868
rect 13142 4924 13206 4928
rect 13142 4868 13146 4924
rect 13146 4868 13202 4924
rect 13202 4868 13206 4924
rect 13142 4864 13206 4868
rect 13222 4924 13286 4928
rect 13222 4868 13226 4924
rect 13226 4868 13282 4924
rect 13282 4868 13286 4924
rect 13222 4864 13286 4868
rect 13302 4924 13366 4928
rect 13302 4868 13306 4924
rect 13306 4868 13362 4924
rect 13362 4868 13366 4924
rect 13302 4864 13366 4868
rect 13382 4924 13446 4928
rect 13382 4868 13386 4924
rect 13386 4868 13442 4924
rect 13442 4868 13446 4924
rect 13382 4864 13446 4868
rect 5828 4380 5892 4384
rect 5828 4324 5832 4380
rect 5832 4324 5888 4380
rect 5888 4324 5892 4380
rect 5828 4320 5892 4324
rect 5908 4380 5972 4384
rect 5908 4324 5912 4380
rect 5912 4324 5968 4380
rect 5968 4324 5972 4380
rect 5908 4320 5972 4324
rect 5988 4380 6052 4384
rect 5988 4324 5992 4380
rect 5992 4324 6048 4380
rect 6048 4324 6052 4380
rect 5988 4320 6052 4324
rect 6068 4380 6132 4384
rect 6068 4324 6072 4380
rect 6072 4324 6128 4380
rect 6128 4324 6132 4380
rect 6068 4320 6132 4324
rect 10704 4380 10768 4384
rect 10704 4324 10708 4380
rect 10708 4324 10764 4380
rect 10764 4324 10768 4380
rect 10704 4320 10768 4324
rect 10784 4380 10848 4384
rect 10784 4324 10788 4380
rect 10788 4324 10844 4380
rect 10844 4324 10848 4380
rect 10784 4320 10848 4324
rect 10864 4380 10928 4384
rect 10864 4324 10868 4380
rect 10868 4324 10924 4380
rect 10924 4324 10928 4380
rect 10864 4320 10928 4324
rect 10944 4380 11008 4384
rect 10944 4324 10948 4380
rect 10948 4324 11004 4380
rect 11004 4324 11008 4380
rect 10944 4320 11008 4324
rect 3390 3836 3454 3840
rect 3390 3780 3394 3836
rect 3394 3780 3450 3836
rect 3450 3780 3454 3836
rect 3390 3776 3454 3780
rect 3470 3836 3534 3840
rect 3470 3780 3474 3836
rect 3474 3780 3530 3836
rect 3530 3780 3534 3836
rect 3470 3776 3534 3780
rect 3550 3836 3614 3840
rect 3550 3780 3554 3836
rect 3554 3780 3610 3836
rect 3610 3780 3614 3836
rect 3550 3776 3614 3780
rect 3630 3836 3694 3840
rect 3630 3780 3634 3836
rect 3634 3780 3690 3836
rect 3690 3780 3694 3836
rect 3630 3776 3694 3780
rect 8266 3836 8330 3840
rect 8266 3780 8270 3836
rect 8270 3780 8326 3836
rect 8326 3780 8330 3836
rect 8266 3776 8330 3780
rect 8346 3836 8410 3840
rect 8346 3780 8350 3836
rect 8350 3780 8406 3836
rect 8406 3780 8410 3836
rect 8346 3776 8410 3780
rect 8426 3836 8490 3840
rect 8426 3780 8430 3836
rect 8430 3780 8486 3836
rect 8486 3780 8490 3836
rect 8426 3776 8490 3780
rect 8506 3836 8570 3840
rect 8506 3780 8510 3836
rect 8510 3780 8566 3836
rect 8566 3780 8570 3836
rect 8506 3776 8570 3780
rect 13142 3836 13206 3840
rect 13142 3780 13146 3836
rect 13146 3780 13202 3836
rect 13202 3780 13206 3836
rect 13142 3776 13206 3780
rect 13222 3836 13286 3840
rect 13222 3780 13226 3836
rect 13226 3780 13282 3836
rect 13282 3780 13286 3836
rect 13222 3776 13286 3780
rect 13302 3836 13366 3840
rect 13302 3780 13306 3836
rect 13306 3780 13362 3836
rect 13362 3780 13366 3836
rect 13302 3776 13366 3780
rect 13382 3836 13446 3840
rect 13382 3780 13386 3836
rect 13386 3780 13442 3836
rect 13442 3780 13446 3836
rect 13382 3776 13446 3780
rect 5828 3292 5892 3296
rect 5828 3236 5832 3292
rect 5832 3236 5888 3292
rect 5888 3236 5892 3292
rect 5828 3232 5892 3236
rect 5908 3292 5972 3296
rect 5908 3236 5912 3292
rect 5912 3236 5968 3292
rect 5968 3236 5972 3292
rect 5908 3232 5972 3236
rect 5988 3292 6052 3296
rect 5988 3236 5992 3292
rect 5992 3236 6048 3292
rect 6048 3236 6052 3292
rect 5988 3232 6052 3236
rect 6068 3292 6132 3296
rect 6068 3236 6072 3292
rect 6072 3236 6128 3292
rect 6128 3236 6132 3292
rect 6068 3232 6132 3236
rect 10704 3292 10768 3296
rect 10704 3236 10708 3292
rect 10708 3236 10764 3292
rect 10764 3236 10768 3292
rect 10704 3232 10768 3236
rect 10784 3292 10848 3296
rect 10784 3236 10788 3292
rect 10788 3236 10844 3292
rect 10844 3236 10848 3292
rect 10784 3232 10848 3236
rect 10864 3292 10928 3296
rect 10864 3236 10868 3292
rect 10868 3236 10924 3292
rect 10924 3236 10928 3292
rect 10864 3232 10928 3236
rect 10944 3292 11008 3296
rect 10944 3236 10948 3292
rect 10948 3236 11004 3292
rect 11004 3236 11008 3292
rect 10944 3232 11008 3236
rect 3390 2748 3454 2752
rect 3390 2692 3394 2748
rect 3394 2692 3450 2748
rect 3450 2692 3454 2748
rect 3390 2688 3454 2692
rect 3470 2748 3534 2752
rect 3470 2692 3474 2748
rect 3474 2692 3530 2748
rect 3530 2692 3534 2748
rect 3470 2688 3534 2692
rect 3550 2748 3614 2752
rect 3550 2692 3554 2748
rect 3554 2692 3610 2748
rect 3610 2692 3614 2748
rect 3550 2688 3614 2692
rect 3630 2748 3694 2752
rect 3630 2692 3634 2748
rect 3634 2692 3690 2748
rect 3690 2692 3694 2748
rect 3630 2688 3694 2692
rect 8266 2748 8330 2752
rect 8266 2692 8270 2748
rect 8270 2692 8326 2748
rect 8326 2692 8330 2748
rect 8266 2688 8330 2692
rect 8346 2748 8410 2752
rect 8346 2692 8350 2748
rect 8350 2692 8406 2748
rect 8406 2692 8410 2748
rect 8346 2688 8410 2692
rect 8426 2748 8490 2752
rect 8426 2692 8430 2748
rect 8430 2692 8486 2748
rect 8486 2692 8490 2748
rect 8426 2688 8490 2692
rect 8506 2748 8570 2752
rect 8506 2692 8510 2748
rect 8510 2692 8566 2748
rect 8566 2692 8570 2748
rect 8506 2688 8570 2692
rect 13142 2748 13206 2752
rect 13142 2692 13146 2748
rect 13146 2692 13202 2748
rect 13202 2692 13206 2748
rect 13142 2688 13206 2692
rect 13222 2748 13286 2752
rect 13222 2692 13226 2748
rect 13226 2692 13282 2748
rect 13282 2692 13286 2748
rect 13222 2688 13286 2692
rect 13302 2748 13366 2752
rect 13302 2692 13306 2748
rect 13306 2692 13362 2748
rect 13362 2692 13366 2748
rect 13302 2688 13366 2692
rect 13382 2748 13446 2752
rect 13382 2692 13386 2748
rect 13386 2692 13442 2748
rect 13442 2692 13446 2748
rect 13382 2688 13446 2692
rect 5828 2204 5892 2208
rect 5828 2148 5832 2204
rect 5832 2148 5888 2204
rect 5888 2148 5892 2204
rect 5828 2144 5892 2148
rect 5908 2204 5972 2208
rect 5908 2148 5912 2204
rect 5912 2148 5968 2204
rect 5968 2148 5972 2204
rect 5908 2144 5972 2148
rect 5988 2204 6052 2208
rect 5988 2148 5992 2204
rect 5992 2148 6048 2204
rect 6048 2148 6052 2204
rect 5988 2144 6052 2148
rect 6068 2204 6132 2208
rect 6068 2148 6072 2204
rect 6072 2148 6128 2204
rect 6128 2148 6132 2204
rect 6068 2144 6132 2148
rect 10704 2204 10768 2208
rect 10704 2148 10708 2204
rect 10708 2148 10764 2204
rect 10764 2148 10768 2204
rect 10704 2144 10768 2148
rect 10784 2204 10848 2208
rect 10784 2148 10788 2204
rect 10788 2148 10844 2204
rect 10844 2148 10848 2204
rect 10784 2144 10848 2148
rect 10864 2204 10928 2208
rect 10864 2148 10868 2204
rect 10868 2148 10924 2204
rect 10924 2148 10928 2204
rect 10864 2144 10928 2148
rect 10944 2204 11008 2208
rect 10944 2148 10948 2204
rect 10948 2148 11004 2204
rect 11004 2148 11008 2204
rect 10944 2144 11008 2148
<< metal4 >>
rect 3382 15808 3702 16368
rect 3382 15744 3390 15808
rect 3454 15744 3470 15808
rect 3534 15744 3550 15808
rect 3614 15744 3630 15808
rect 3694 15744 3702 15808
rect 3382 14720 3702 15744
rect 3382 14656 3390 14720
rect 3454 14656 3470 14720
rect 3534 14656 3550 14720
rect 3614 14656 3630 14720
rect 3694 14656 3702 14720
rect 3382 14032 3702 14656
rect 3382 13796 3424 14032
rect 3660 13796 3702 14032
rect 3382 13632 3702 13796
rect 3382 13568 3390 13632
rect 3454 13568 3470 13632
rect 3534 13568 3550 13632
rect 3614 13568 3630 13632
rect 3694 13568 3702 13632
rect 3382 12544 3702 13568
rect 3382 12480 3390 12544
rect 3454 12480 3470 12544
rect 3534 12480 3550 12544
rect 3614 12480 3630 12544
rect 3694 12480 3702 12544
rect 3382 11456 3702 12480
rect 3382 11392 3390 11456
rect 3454 11392 3470 11456
rect 3534 11392 3550 11456
rect 3614 11392 3630 11456
rect 3694 11392 3702 11456
rect 3382 10368 3702 11392
rect 3382 10304 3390 10368
rect 3454 10304 3470 10368
rect 3534 10304 3550 10368
rect 3614 10304 3630 10368
rect 3694 10304 3702 10368
rect 3382 9318 3702 10304
rect 3382 9280 3424 9318
rect 3660 9280 3702 9318
rect 3382 9216 3390 9280
rect 3694 9216 3702 9280
rect 3382 9082 3424 9216
rect 3660 9082 3702 9216
rect 3382 8192 3702 9082
rect 3382 8128 3390 8192
rect 3454 8128 3470 8192
rect 3534 8128 3550 8192
rect 3614 8128 3630 8192
rect 3694 8128 3702 8192
rect 3382 7104 3702 8128
rect 3382 7040 3390 7104
rect 3454 7040 3470 7104
rect 3534 7040 3550 7104
rect 3614 7040 3630 7104
rect 3694 7040 3702 7104
rect 3382 6016 3702 7040
rect 3382 5952 3390 6016
rect 3454 5952 3470 6016
rect 3534 5952 3550 6016
rect 3614 5952 3630 6016
rect 3694 5952 3702 6016
rect 3382 4928 3702 5952
rect 3382 4864 3390 4928
rect 3454 4864 3470 4928
rect 3534 4864 3550 4928
rect 3614 4864 3630 4928
rect 3694 4864 3702 4928
rect 3382 4603 3702 4864
rect 3382 4367 3424 4603
rect 3660 4367 3702 4603
rect 3382 3840 3702 4367
rect 3382 3776 3390 3840
rect 3454 3776 3470 3840
rect 3534 3776 3550 3840
rect 3614 3776 3630 3840
rect 3694 3776 3702 3840
rect 3382 2752 3702 3776
rect 3382 2688 3390 2752
rect 3454 2688 3470 2752
rect 3534 2688 3550 2752
rect 3614 2688 3630 2752
rect 3694 2688 3702 2752
rect 3382 2128 3702 2688
rect 5820 16352 6140 16368
rect 5820 16288 5828 16352
rect 5892 16288 5908 16352
rect 5972 16288 5988 16352
rect 6052 16288 6068 16352
rect 6132 16288 6140 16352
rect 5820 15264 6140 16288
rect 5820 15200 5828 15264
rect 5892 15200 5908 15264
rect 5972 15200 5988 15264
rect 6052 15200 6068 15264
rect 6132 15200 6140 15264
rect 5820 14176 6140 15200
rect 5820 14112 5828 14176
rect 5892 14112 5908 14176
rect 5972 14112 5988 14176
rect 6052 14112 6068 14176
rect 6132 14112 6140 14176
rect 5820 13088 6140 14112
rect 5820 13024 5828 13088
rect 5892 13024 5908 13088
rect 5972 13024 5988 13088
rect 6052 13024 6068 13088
rect 6132 13024 6140 13088
rect 5820 12000 6140 13024
rect 5820 11936 5828 12000
rect 5892 11936 5908 12000
rect 5972 11936 5988 12000
rect 6052 11936 6068 12000
rect 6132 11936 6140 12000
rect 5820 11675 6140 11936
rect 5820 11439 5862 11675
rect 6098 11439 6140 11675
rect 5820 10912 6140 11439
rect 5820 10848 5828 10912
rect 5892 10848 5908 10912
rect 5972 10848 5988 10912
rect 6052 10848 6068 10912
rect 6132 10848 6140 10912
rect 5820 9824 6140 10848
rect 5820 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6140 9824
rect 5820 8736 6140 9760
rect 5820 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6140 8736
rect 5820 7648 6140 8672
rect 5820 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6140 7648
rect 5820 6960 6140 7584
rect 5820 6724 5862 6960
rect 6098 6724 6140 6960
rect 5820 6560 6140 6724
rect 5820 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6140 6560
rect 5820 5472 6140 6496
rect 5820 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6140 5472
rect 5820 4384 6140 5408
rect 5820 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6140 4384
rect 5820 3296 6140 4320
rect 5820 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6140 3296
rect 5820 2208 6140 3232
rect 5820 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6140 2208
rect 5820 2128 6140 2144
rect 8258 15808 8578 16368
rect 8258 15744 8266 15808
rect 8330 15744 8346 15808
rect 8410 15744 8426 15808
rect 8490 15744 8506 15808
rect 8570 15744 8578 15808
rect 8258 14720 8578 15744
rect 8258 14656 8266 14720
rect 8330 14656 8346 14720
rect 8410 14656 8426 14720
rect 8490 14656 8506 14720
rect 8570 14656 8578 14720
rect 8258 14032 8578 14656
rect 8258 13796 8300 14032
rect 8536 13796 8578 14032
rect 8258 13632 8578 13796
rect 8258 13568 8266 13632
rect 8330 13568 8346 13632
rect 8410 13568 8426 13632
rect 8490 13568 8506 13632
rect 8570 13568 8578 13632
rect 8258 12544 8578 13568
rect 8258 12480 8266 12544
rect 8330 12480 8346 12544
rect 8410 12480 8426 12544
rect 8490 12480 8506 12544
rect 8570 12480 8578 12544
rect 8258 11456 8578 12480
rect 8258 11392 8266 11456
rect 8330 11392 8346 11456
rect 8410 11392 8426 11456
rect 8490 11392 8506 11456
rect 8570 11392 8578 11456
rect 8258 10368 8578 11392
rect 8258 10304 8266 10368
rect 8330 10304 8346 10368
rect 8410 10304 8426 10368
rect 8490 10304 8506 10368
rect 8570 10304 8578 10368
rect 8258 9318 8578 10304
rect 8258 9280 8300 9318
rect 8536 9280 8578 9318
rect 8258 9216 8266 9280
rect 8570 9216 8578 9280
rect 8258 9082 8300 9216
rect 8536 9082 8578 9216
rect 8258 8192 8578 9082
rect 8258 8128 8266 8192
rect 8330 8128 8346 8192
rect 8410 8128 8426 8192
rect 8490 8128 8506 8192
rect 8570 8128 8578 8192
rect 8258 7104 8578 8128
rect 8258 7040 8266 7104
rect 8330 7040 8346 7104
rect 8410 7040 8426 7104
rect 8490 7040 8506 7104
rect 8570 7040 8578 7104
rect 8258 6016 8578 7040
rect 8258 5952 8266 6016
rect 8330 5952 8346 6016
rect 8410 5952 8426 6016
rect 8490 5952 8506 6016
rect 8570 5952 8578 6016
rect 8258 4928 8578 5952
rect 8258 4864 8266 4928
rect 8330 4864 8346 4928
rect 8410 4864 8426 4928
rect 8490 4864 8506 4928
rect 8570 4864 8578 4928
rect 8258 4603 8578 4864
rect 8258 4367 8300 4603
rect 8536 4367 8578 4603
rect 8258 3840 8578 4367
rect 8258 3776 8266 3840
rect 8330 3776 8346 3840
rect 8410 3776 8426 3840
rect 8490 3776 8506 3840
rect 8570 3776 8578 3840
rect 8258 2752 8578 3776
rect 8258 2688 8266 2752
rect 8330 2688 8346 2752
rect 8410 2688 8426 2752
rect 8490 2688 8506 2752
rect 8570 2688 8578 2752
rect 8258 2128 8578 2688
rect 10696 16352 11016 16368
rect 10696 16288 10704 16352
rect 10768 16288 10784 16352
rect 10848 16288 10864 16352
rect 10928 16288 10944 16352
rect 11008 16288 11016 16352
rect 10696 15264 11016 16288
rect 10696 15200 10704 15264
rect 10768 15200 10784 15264
rect 10848 15200 10864 15264
rect 10928 15200 10944 15264
rect 11008 15200 11016 15264
rect 10696 14176 11016 15200
rect 10696 14112 10704 14176
rect 10768 14112 10784 14176
rect 10848 14112 10864 14176
rect 10928 14112 10944 14176
rect 11008 14112 11016 14176
rect 10696 13088 11016 14112
rect 10696 13024 10704 13088
rect 10768 13024 10784 13088
rect 10848 13024 10864 13088
rect 10928 13024 10944 13088
rect 11008 13024 11016 13088
rect 10696 12000 11016 13024
rect 10696 11936 10704 12000
rect 10768 11936 10784 12000
rect 10848 11936 10864 12000
rect 10928 11936 10944 12000
rect 11008 11936 11016 12000
rect 10696 11675 11016 11936
rect 10696 11439 10738 11675
rect 10974 11439 11016 11675
rect 10696 10912 11016 11439
rect 10696 10848 10704 10912
rect 10768 10848 10784 10912
rect 10848 10848 10864 10912
rect 10928 10848 10944 10912
rect 11008 10848 11016 10912
rect 10696 9824 11016 10848
rect 10696 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11016 9824
rect 10696 8736 11016 9760
rect 10696 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11016 8736
rect 10696 7648 11016 8672
rect 10696 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11016 7648
rect 10696 6960 11016 7584
rect 10696 6724 10738 6960
rect 10974 6724 11016 6960
rect 10696 6560 11016 6724
rect 10696 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11016 6560
rect 10696 5472 11016 6496
rect 10696 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11016 5472
rect 10696 4384 11016 5408
rect 10696 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11016 4384
rect 10696 3296 11016 4320
rect 10696 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11016 3296
rect 10696 2208 11016 3232
rect 10696 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11016 2208
rect 10696 2128 11016 2144
rect 13134 15808 13454 16368
rect 13134 15744 13142 15808
rect 13206 15744 13222 15808
rect 13286 15744 13302 15808
rect 13366 15744 13382 15808
rect 13446 15744 13454 15808
rect 13134 14720 13454 15744
rect 13134 14656 13142 14720
rect 13206 14656 13222 14720
rect 13286 14656 13302 14720
rect 13366 14656 13382 14720
rect 13446 14656 13454 14720
rect 13134 14032 13454 14656
rect 13134 13796 13176 14032
rect 13412 13796 13454 14032
rect 13134 13632 13454 13796
rect 13134 13568 13142 13632
rect 13206 13568 13222 13632
rect 13286 13568 13302 13632
rect 13366 13568 13382 13632
rect 13446 13568 13454 13632
rect 13134 12544 13454 13568
rect 13134 12480 13142 12544
rect 13206 12480 13222 12544
rect 13286 12480 13302 12544
rect 13366 12480 13382 12544
rect 13446 12480 13454 12544
rect 13134 11456 13454 12480
rect 13134 11392 13142 11456
rect 13206 11392 13222 11456
rect 13286 11392 13302 11456
rect 13366 11392 13382 11456
rect 13446 11392 13454 11456
rect 13134 10368 13454 11392
rect 13134 10304 13142 10368
rect 13206 10304 13222 10368
rect 13286 10304 13302 10368
rect 13366 10304 13382 10368
rect 13446 10304 13454 10368
rect 13134 9318 13454 10304
rect 13134 9280 13176 9318
rect 13412 9280 13454 9318
rect 13134 9216 13142 9280
rect 13446 9216 13454 9280
rect 13134 9082 13176 9216
rect 13412 9082 13454 9216
rect 13134 8192 13454 9082
rect 13134 8128 13142 8192
rect 13206 8128 13222 8192
rect 13286 8128 13302 8192
rect 13366 8128 13382 8192
rect 13446 8128 13454 8192
rect 13134 7104 13454 8128
rect 13134 7040 13142 7104
rect 13206 7040 13222 7104
rect 13286 7040 13302 7104
rect 13366 7040 13382 7104
rect 13446 7040 13454 7104
rect 13134 6016 13454 7040
rect 13134 5952 13142 6016
rect 13206 5952 13222 6016
rect 13286 5952 13302 6016
rect 13366 5952 13382 6016
rect 13446 5952 13454 6016
rect 13134 4928 13454 5952
rect 13134 4864 13142 4928
rect 13206 4864 13222 4928
rect 13286 4864 13302 4928
rect 13366 4864 13382 4928
rect 13446 4864 13454 4928
rect 13134 4603 13454 4864
rect 13134 4367 13176 4603
rect 13412 4367 13454 4603
rect 13134 3840 13454 4367
rect 13134 3776 13142 3840
rect 13206 3776 13222 3840
rect 13286 3776 13302 3840
rect 13366 3776 13382 3840
rect 13446 3776 13454 3840
rect 13134 2752 13454 3776
rect 13134 2688 13142 2752
rect 13206 2688 13222 2752
rect 13286 2688 13302 2752
rect 13366 2688 13382 2752
rect 13446 2688 13454 2752
rect 13134 2128 13454 2688
<< via4 >>
rect 3424 13796 3660 14032
rect 3424 9280 3660 9318
rect 3424 9216 3454 9280
rect 3454 9216 3470 9280
rect 3470 9216 3534 9280
rect 3534 9216 3550 9280
rect 3550 9216 3614 9280
rect 3614 9216 3630 9280
rect 3630 9216 3660 9280
rect 3424 9082 3660 9216
rect 3424 4367 3660 4603
rect 5862 11439 6098 11675
rect 5862 6724 6098 6960
rect 8300 13796 8536 14032
rect 8300 9280 8536 9318
rect 8300 9216 8330 9280
rect 8330 9216 8346 9280
rect 8346 9216 8410 9280
rect 8410 9216 8426 9280
rect 8426 9216 8490 9280
rect 8490 9216 8506 9280
rect 8506 9216 8536 9280
rect 8300 9082 8536 9216
rect 8300 4367 8536 4603
rect 10738 11439 10974 11675
rect 10738 6724 10974 6960
rect 13176 13796 13412 14032
rect 13176 9280 13412 9318
rect 13176 9216 13206 9280
rect 13206 9216 13222 9280
rect 13222 9216 13286 9280
rect 13286 9216 13302 9280
rect 13302 9216 13366 9280
rect 13366 9216 13382 9280
rect 13382 9216 13412 9280
rect 13176 9082 13412 9216
rect 13176 4367 13412 4603
<< metal5 >>
rect 1104 14032 15732 14074
rect 1104 13796 3424 14032
rect 3660 13796 8300 14032
rect 8536 13796 13176 14032
rect 13412 13796 15732 14032
rect 1104 13754 15732 13796
rect 1104 11675 15732 11717
rect 1104 11439 5862 11675
rect 6098 11439 10738 11675
rect 10974 11439 15732 11675
rect 1104 11397 15732 11439
rect 1104 9318 15732 9360
rect 1104 9082 3424 9318
rect 3660 9082 8300 9318
rect 8536 9082 13176 9318
rect 13412 9082 15732 9318
rect 1104 9040 15732 9082
rect 1104 6960 15732 7002
rect 1104 6724 5862 6960
rect 6098 6724 10738 6960
rect 10974 6724 15732 6960
rect 1104 6682 15732 6724
rect 1104 4603 15732 4646
rect 1104 4367 3424 4603
rect 3660 4367 8300 4603
rect 8536 4367 13176 4603
rect 13412 4367 15732 4603
rect 1104 4325 15732 4367
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1629722742
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1629722742
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1629722742
transform 1 0 1380 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1629722742
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1629722742
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1629722742
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1629722742
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1629722742
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _434_
timestamp 1629722742
transform -1 0 4048 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _453_
timestamp 1629722742
transform 1 0 2668 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output20
timestamp 1629722742
transform -1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36
timestamp 1629722742
transform 1 0 4416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_32
timestamp 1629722742
transform 1 0 4048 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1629722742
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _454_
timestamp 1629722742
transform -1 0 4416 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output21
timestamp 1629722742
transform -1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47
timestamp 1629722742
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1629722742
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_44
timestamp 1629722742
transform 1 0 5152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _452_
timestamp 1629722742
transform -1 0 5888 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2oi_1  _467_
timestamp 1629722742
transform -1 0 5428 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1629722742
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1629722742
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1629722742
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1629722742
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1629722742
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1629722742
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1629722742
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_63
timestamp 1629722742
transform 1 0 6900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output24
timestamp 1629722742
transform -1 0 6900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _431_
timestamp 1629722742
transform 1 0 6808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70
timestamp 1629722742
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77
timestamp 1629722742
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1629722742
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _428_
timestamp 1629722742
transform -1 0 8004 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1629722742
transform 1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1629722742
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_79
timestamp 1629722742
transform 1 0 8372 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_84
timestamp 1629722742
transform 1 0 8832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1629722742
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _445_
timestamp 1629722742
transform 1 0 9200 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _447_
timestamp 1629722742
transform -1 0 8832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _449_
timestamp 1629722742
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101
timestamp 1629722742
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93
timestamp 1629722742
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1629722742
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _427_
timestamp 1629722742
transform 1 0 10304 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output29
timestamp 1629722742
transform -1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1629722742
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1629722742
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1629722742
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1629722742
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1629722742
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _438_
timestamp 1629722742
transform -1 0 12144 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1629722742
transform -1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1629722742
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128
timestamp 1629722742
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_116
timestamp 1629722742
transform 1 0 11776 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2ai_2  _465_
timestamp 1629722742
transform -1 0 13248 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output19
timestamp 1629722742
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1629722742
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 1629722742
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1629722742
transform 1 0 13248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1629722742
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_2  _473_
timestamp 1629722742
transform -1 0 14720 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1629722742
transform -1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152
timestamp 1629722742
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_148
timestamp 1629722742
transform 1 0 14720 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _471_
timestamp 1629722742
transform -1 0 15088 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1629722742
transform -1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1629722742
transform -1 0 15732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1629722742
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1629722742
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1629722742
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _436_
timestamp 1629722742
transform 1 0 1840 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_2_15
timestamp 1629722742
transform 1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1629722742
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1629722742
transform -1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_32
timestamp 1629722742
transform 1 0 4048 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1629722742
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1629722742
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _466_
timestamp 1629722742
transform 1 0 4600 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_2_45
timestamp 1629722742
transform 1 0 5244 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_53
timestamp 1629722742
transform 1 0 5980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1629722742
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _420_
timestamp 1629722742
transform 1 0 6164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _437_
timestamp 1629722742
transform 1 0 6808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1629722742
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1629722742
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _430_
timestamp 1629722742
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1629722742
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1629722742
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1629722742
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _455_
timestamp 1629722742
transform -1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_97
timestamp 1629722742
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_105
timestamp 1629722742
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_113
timestamp 1629722742
transform 1 0 11500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _426_
timestamp 1629722742
transform 1 0 10856 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_2_124
timestamp 1629722742
transform 1 0 12512 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _472_
timestamp 1629722742
transform -1 0 12512 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1629722742
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1629722742
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _474_
timestamp 1629722742
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output23
timestamp 1629722742
transform 1 0 13248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_149
timestamp 1629722742
transform 1 0 14812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_155
timestamp 1629722742
transform 1 0 15364 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1629722742
transform -1 0 15732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1629722742
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1629722742
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1629722742
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _435_
timestamp 1629722742
transform 1 0 1840 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_3_15
timestamp 1629722742
transform 1 0 2484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1629722742
transform 1 0 3312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1629722742
transform -1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_36
timestamp 1629722742
transform 1 0 4416 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _415_
timestamp 1629722742
transform 1 0 3680 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _413_
timestamp 1629722742
transform 1 0 5152 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1629722742
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_60
timestamp 1629722742
transform 1 0 6624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1629722742
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1629722742
transform -1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _421_
timestamp 1629722742
transform -1 0 7636 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_3_71
timestamp 1629722742
transform 1 0 7636 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _448_
timestamp 1629722742
transform -1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_80
timestamp 1629722742
transform 1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_87
timestamp 1629722742
transform 1 0 9108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _399_
timestamp 1629722742
transform -1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_101
timestamp 1629722742
transform 1 0 10396 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp 1629722742
transform 1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 1629722742
transform 1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1629722742
transform 1 0 9476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1629722742
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1629722742
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1629722742
transform -1 0 11040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _409_
timestamp 1629722742
transform -1 0 12144 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_3_120
timestamp 1629722742
transform 1 0 12144 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _463_
timestamp 1629722742
transform 1 0 12880 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_3_133
timestamp 1629722742
transform 1 0 13340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_137
timestamp 1629722742
transform 1 0 13708 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _468_
timestamp 1629722742
transform -1 0 14536 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_146
timestamp 1629722742
transform 1 0 14536 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_154
timestamp 1629722742
transform 1 0 15272 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1629722742
transform -1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1629722742
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1629722742
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _418_
timestamp 1629722742
transform 1 0 1380 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_4_14
timestamp 1629722742
transform 1 0 2392 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_22
timestamp 1629722742
transform 1 0 3128 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2ai_1  _416_
timestamp 1629722742
transform -1 0 3128 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1629722742
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1629722742
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _414_
timestamp 1629722742
transform 1 0 4140 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1629722742
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _401_
timestamp 1629722742
transform 1 0 5244 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1629722742
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_60
timestamp 1629722742
transform 1 0 6624 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_64
timestamp 1629722742
transform 1 0 6992 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _400_
timestamp 1629722742
transform 1 0 6348 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_73
timestamp 1629722742
transform 1 0 7820 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _369_
timestamp 1629722742
transform -1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _412_
timestamp 1629722742
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1629722742
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp 1629722742
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1629722742
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _424_
timestamp 1629722742
transform -1 0 9844 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_4_95
timestamp 1629722742
transform 1 0 9844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _379_
timestamp 1629722742
transform -1 0 10672 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_4_104
timestamp 1629722742
transform 1 0 10672 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _422_
timestamp 1629722742
transform 1 0 11224 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_118
timestamp 1629722742
transform 1 0 11960 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1629722742
transform 1 0 12696 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_1  _464_
timestamp 1629722742
transform 1 0 12880 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1629722742
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1629722742
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1629722742
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_151
timestamp 1629722742
transform 1 0 14996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _461_
timestamp 1629722742
transform -1 0 14996 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_155
timestamp 1629722742
transform 1 0 15364 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1629722742
transform -1 0 15732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_6
timestamp 1629722742
transform 1 0 1656 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1629722742
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1629722742
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_17
timestamp 1629722742
transform 1 0 2668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1629722742
transform 1 0 3312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _502_
timestamp 1629722742
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1629722742
transform 1 0 2392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_35
timestamp 1629722742
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _419_
timestamp 1629722742
transform 1 0 3680 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_5_46
timestamp 1629722742
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _402_
timestamp 1629722742
transform 1 0 4692 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1629722742
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 1629722742
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1629722742
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _372_
timestamp 1629722742
transform 1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_66
timestamp 1629722742
transform 1 0 7176 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _370_
timestamp 1629722742
transform 1 0 7728 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_5_79
timestamp 1629722742
transform 1 0 8372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _397_
timestamp 1629722742
transform -1 0 9384 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_5_90
timestamp 1629722742
transform 1 0 9384 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _381_
timestamp 1629722742
transform -1 0 10580 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1629722742
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1629722742
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1629722742
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1629722742
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _406_
timestamp 1629722742
transform 1 0 11592 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_5_121
timestamp 1629722742
transform 1 0 12236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _443_
timestamp 1629722742
transform 1 0 12788 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_5_132
timestamp 1629722742
transform 1 0 13248 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_140
timestamp 1629722742
transform 1 0 13984 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _439_
timestamp 1629722742
transform 1 0 14076 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_144
timestamp 1629722742
transform 1 0 14352 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_152
timestamp 1629722742
transform 1 0 15088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output32
timestamp 1629722742
transform 1 0 14720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1629722742
transform -1 0 15732 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_10
timestamp 1629722742
transform 1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1629722742
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1629722742
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1629722742
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _395_
timestamp 1629722742
transform -1 0 2392 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _417_
timestamp 1629722742
transform 1 0 1380 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1629722742
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1629722742
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_14
timestamp 1629722742
transform 1 0 2392 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_22
timestamp 1629722742
transform 1 0 3128 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_1  _391_
timestamp 1629722742
transform -1 0 4048 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1629722742
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1629722742
transform 1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_37
timestamp 1629722742
transform 1 0 4508 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_32
timestamp 1629722742
transform 1 0 4048 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1629722742
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _390_
timestamp 1629722742
transform 1 0 4416 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _392_
timestamp 1629722742
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_46
timestamp 1629722742
transform 1 0 5336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_44
timestamp 1629722742
transform 1 0 5152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_48
timestamp 1629722742
transform 1 0 5520 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _373_
timestamp 1629722742
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _374_
timestamp 1629722742
transform 1 0 5704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1629722742
transform -1 0 5336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1629722742
transform 1 0 6440 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1629722742
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1629722742
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1629722742
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__and4_1  _371_
timestamp 1629722742
transform -1 0 7360 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _411_
timestamp 1629722742
transform -1 0 7176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_66
timestamp 1629722742
transform 1 0 7176 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_72
timestamp 1629722742
transform 1 0 7728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_68
timestamp 1629722742
transform 1 0 7360 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _386_
timestamp 1629722742
transform 1 0 7912 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _410_
timestamp 1629722742
transform 1 0 7820 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1629722742
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1629722742
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_82
timestamp 1629722742
transform 1 0 8648 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_88
timestamp 1629722742
transform 1 0 9200 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1629722742
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _383_
timestamp 1629722742
transform -1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _398_
timestamp 1629722742
transform -1 0 9936 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_101
timestamp 1629722742
transform 1 0 10396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1629722742
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_102
timestamp 1629722742
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_96
timestamp 1629722742
transform 1 0 9936 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _380_
timestamp 1629722742
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_108
timestamp 1629722742
transform 1 0 11040 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_115
timestamp 1629722742
transform 1 0 11684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1629722742
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1629722742
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1629722742
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _377_
timestamp 1629722742
transform -1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _382_
timestamp 1629722742
transform 1 0 11408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _403_
timestamp 1629722742
transform 1 0 10580 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _405_
timestamp 1629722742
transform -1 0 12236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_122
timestamp 1629722742
transform 1 0 12328 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_121
timestamp 1629722742
transform 1 0 12236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _404_
timestamp 1629722742
transform 1 0 12052 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1629722742
transform -1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _444_
timestamp 1629722742
transform 1 0 12604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_129
timestamp 1629722742
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1629722742
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 1629722742
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1629722742
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_137
timestamp 1629722742
transform 1 0 13708 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1629722742
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 1629722742
transform -1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _458_
timestamp 1629722742
transform -1 0 14536 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_150
timestamp 1629722742
transform 1 0 14904 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_146
timestamp 1629722742
transform 1 0 14536 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_154
timestamp 1629722742
transform 1 0 15272 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_1  _440_
timestamp 1629722742
transform -1 0 14904 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1629722742
transform -1 0 15732 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1629722742
transform -1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1629722742
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1629722742
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1629722742
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _393_
timestamp 1629722742
transform -1 0 2484 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1629722742
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1629722742
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_36
timestamp 1629722742
transform 1 0 4416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1629722742
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _396_
timestamp 1629722742
transform 1 0 3772 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_8_40
timestamp 1629722742
transform 1 0 4784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_49
timestamp 1629722742
transform 1 0 5612 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _389_
timestamp 1629722742
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_63
timestamp 1629722742
transform 1 0 6900 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _388_
timestamp 1629722742
transform 1 0 6164 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_69
timestamp 1629722742
transform 1 0 7452 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_73
timestamp 1629722742
transform 1 0 7820 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _347_
timestamp 1629722742
transform 1 0 7544 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _460_
timestamp 1629722742
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1629722742
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1629722742
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _385_
timestamp 1629722742
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1629722742
transform 1 0 9660 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_97
timestamp 1629722742
transform 1 0 10028 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _344_
timestamp 1629722742
transform 1 0 10120 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_8_103
timestamp 1629722742
transform 1 0 10580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_115
timestamp 1629722742
transform 1 0 11684 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _345_
timestamp 1629722742
transform 1 0 10948 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_126
timestamp 1629722742
transform 1 0 12696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _384_
timestamp 1629722742
transform 1 0 12052 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1629722742
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1629722742
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1629722742
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1629722742
transform 1 0 13064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _378_
timestamp 1629722742
transform 1 0 14076 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_8_151
timestamp 1629722742
transform 1 0 14996 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_155
timestamp 1629722742
transform 1 0 15364 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1629722742
transform -1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1629722742
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1629722742
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1629722742
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_22
timestamp 1629722742
transform 1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _527_
timestamp 1629722742
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_33
timestamp 1629722742
transform 1 0 4140 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _375_
timestamp 1629722742
transform 1 0 3496 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_9_41
timestamp 1629722742
transform 1 0 4876 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_50
timestamp 1629722742
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _387_
timestamp 1629722742
transform 1 0 5060 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_9_57
timestamp 1629722742
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1629722742
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _348_
timestamp 1629722742
transform 1 0 6900 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_71
timestamp 1629722742
transform 1 0 7636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1629722742
transform -1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_78
timestamp 1629722742
transform 1 0 8280 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_84
timestamp 1629722742
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_88
timestamp 1629722742
transform 1 0 9200 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1629722742
transform -1 0 9200 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1629722742
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _376_
timestamp 1629722742
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _503_
timestamp 1629722742
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1629722742
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1629722742
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1629722742
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1629722742
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _456_
timestamp 1629722742
transform 1 0 11592 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_117
timestamp 1629722742
transform 1 0 11868 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _343_
timestamp 1629722742
transform 1 0 12236 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_129
timestamp 1629722742
transform 1 0 12972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_136
timestamp 1629722742
transform 1 0 13616 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1629722742
transform 1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _441_
timestamp 1629722742
transform 1 0 13984 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_9_147
timestamp 1629722742
transform 1 0 14628 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_155
timestamp 1629722742
transform 1 0 15364 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1629722742
transform -1 0 15732 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_12
timestamp 1629722742
transform 1 0 2208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1629722742
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1629722742
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _367_
timestamp 1629722742
transform 1 0 1564 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1629722742
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _362_
timestamp 1629722742
transform 1 0 2576 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1629722742
transform 1 0 4048 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1629722742
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _358_
timestamp 1629722742
transform 1 0 4416 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _524_
timestamp 1629722742
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_44
timestamp 1629722742
transform 1 0 5152 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1629722742
transform 1 0 5888 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_62
timestamp 1629722742
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _351_
timestamp 1629722742
transform 1 0 6072 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_69
timestamp 1629722742
transform 1 0 7452 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _339_
timestamp 1629722742
transform -1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1629722742
transform 1 0 7176 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1629722742
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1629722742
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1629722742
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  _356_
timestamp 1629722742
transform 1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_102
timestamp 1629722742
transform 1 0 10488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_93
timestamp 1629722742
transform 1 0 9660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1629722742
transform -1 0 10488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_113
timestamp 1629722742
transform 1 0 11500 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _322_
timestamp 1629722742
transform 1 0 10856 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_10_117
timestamp 1629722742
transform 1 0 11868 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp 1629722742
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _319_
timestamp 1629722742
transform 1 0 11960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _323_
timestamp 1629722742
transform -1 0 13248 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_10_132
timestamp 1629722742
transform 1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1629722742
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1629722742
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_152
timestamp 1629722742
transform 1 0 15088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _321_
timestamp 1629722742
transform 1 0 14168 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1629722742
transform -1 0 15732 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1629722742
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1629722742
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _363_
timestamp 1629722742
transform 1 0 1748 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1629722742
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_23
timestamp 1629722742
transform 1 0 3220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output17
timestamp 1629722742
transform -1 0 3220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_35
timestamp 1629722742
transform 1 0 4324 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _361_
timestamp 1629722742
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_43
timestamp 1629722742
transform 1 0 5060 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _357_
timestamp 1629722742
transform 1 0 5152 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1629722742
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1629722742
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_61
timestamp 1629722742
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1629722742
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _506_
timestamp 1629722742
transform 1 0 6440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_71
timestamp 1629722742
transform 1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _355_
timestamp 1629722742
transform -1 0 7636 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _368_
timestamp 1629722742
transform -1 0 8924 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1629722742
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _326_
timestamp 1629722742
transform 1 0 9292 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_97
timestamp 1629722742
transform 1 0 10028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _324_
timestamp 1629722742
transform 1 0 10396 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_104
timestamp 1629722742
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1629722742
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _294_
timestamp 1629722742
transform 1 0 11500 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_11_120
timestamp 1629722742
transform 1 0 12144 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _342_
timestamp 1629722742
transform -1 0 13340 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_11_133
timestamp 1629722742
transform 1 0 13340 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 1629722742
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _532_
timestamp 1629722742
transform 1 0 13708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_149
timestamp 1629722742
transform 1 0 14812 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _529_
timestamp 1629722742
transform -1 0 14812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_155
timestamp 1629722742
transform 1 0 15364 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1629722742
transform -1 0 15732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1629722742
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1629722742
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _364_
timestamp 1629722742
transform -1 0 2392 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_14
timestamp 1629722742
transform 1 0 2392 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_20
timestamp 1629722742
transform 1 0 2944 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1629722742
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1629722742
transform 1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1629722742
transform 1 0 4048 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1629722742
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _359_
timestamp 1629722742
transform 1 0 4416 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _523_
timestamp 1629722742
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_43
timestamp 1629722742
transform 1 0 5060 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_51
timestamp 1629722742
transform 1 0 5796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_59
timestamp 1629722742
transform 1 0 6532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _318_
timestamp 1629722742
transform -1 0 6532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_67
timestamp 1629722742
transform 1 0 7268 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_75
timestamp 1629722742
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _353_
timestamp 1629722742
transform 1 0 7360 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1629722742
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1629722742
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _293_
timestamp 1629722742
transform 1 0 8924 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_12_90
timestamp 1629722742
transform 1 0 9384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_97
timestamp 1629722742
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _325_
timestamp 1629722742
transform 1 0 9752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_105
timestamp 1629722742
transform 1 0 10764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1629722742
transform 1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _340_
timestamp 1629722742
transform 1 0 11592 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1629722742
transform -1 0 11224 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_119
timestamp 1629722742
transform 1 0 12052 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_125
timestamp 1629722742
transform 1 0 12604 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _485_
timestamp 1629722742
transform -1 0 13156 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_12_131
timestamp 1629722742
transform 1 0 13156 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1629722742
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1629722742
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _528_
timestamp 1629722742
transform 1 0 14076 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_12_146
timestamp 1629722742
transform 1 0 14536 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_154
timestamp 1629722742
transform 1 0 15272 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1629722742
transform -1 0 15732 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1629722742
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1629722742
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp 1629722742
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1629722742
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1629722742
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1629722742
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _297_
timestamp 1629722742
transform 1 0 2024 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output30
timestamp 1629722742
transform -1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_18
timestamp 1629722742
transform 1 0 2760 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1629722742
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _298_
timestamp 1629722742
transform -1 0 3220 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_26
timestamp 1629722742
transform 1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_37
timestamp 1629722742
transform 1 0 4508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1629722742
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1629722742
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_34
timestamp 1629722742
transform 1 0 4232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1629722742
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nand2b_1  _296_
timestamp 1629722742
transform -1 0 5060 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _328_
timestamp 1629722742
transform 1 0 3772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _534_
timestamp 1629722742
transform -1 0 4232 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_49
timestamp 1629722742
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_43
timestamp 1629722742
transform 1 0 5060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_47
timestamp 1629722742
transform 1 0 5428 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_51
timestamp 1629722742
transform 1 0 5796 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _327_
timestamp 1629722742
transform 1 0 4876 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _491_
timestamp 1629722742
transform 1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1629722742
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1629722742
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_55
timestamp 1629722742
transform 1 0 6164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_61
timestamp 1629722742
transform 1 0 6716 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1629722742
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _291_
timestamp 1629722742
transform -1 0 6716 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _316_
timestamp 1629722742
transform 1 0 6624 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_13_67
timestamp 1629722742
transform 1 0 7268 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_71
timestamp 1629722742
transform 1 0 7636 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_69
timestamp 1629722742
transform 1 0 7452 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1629722742
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _290_
timestamp 1629722742
transform 1 0 7728 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _317_
timestamp 1629722742
transform -1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_82
timestamp 1629722742
transform 1 0 8648 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1629722742
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1629722742
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1629722742
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o21ba_1  _299_
timestamp 1629722742
transform 1 0 9108 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_90
timestamp 1629722742
transform 1 0 9384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_98
timestamp 1629722742
transform 1 0 10120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_95
timestamp 1629722742
transform 1 0 9844 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _272_
timestamp 1629722742
transform -1 0 10120 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _496_
timestamp 1629722742
transform 1 0 10488 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1629722742
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1629722742
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_103
timestamp 1629722742
transform 1 0 10580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_112
timestamp 1629722742
transform 1 0 11408 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1629722742
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _271_
timestamp 1629722742
transform 1 0 10764 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _295_
timestamp 1629722742
transform -1 0 12144 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_13_120
timestamp 1629722742
transform 1 0 12144 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_124
timestamp 1629722742
transform 1 0 12512 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_125
timestamp 1629722742
transform 1 0 12604 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _486_
timestamp 1629722742
transform -1 0 13432 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _535_
timestamp 1629722742
transform 1 0 11960 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_13_134
timestamp 1629722742
transform 1 0 13432 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1629722742
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1629722742
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _536_
timestamp 1629722742
transform 1 0 12972 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _547_
timestamp 1629722742
transform 1 0 14076 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_13_142
timestamp 1629722742
transform 1 0 14168 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_151
timestamp 1629722742
transform 1 0 14996 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_151
timestamp 1629722742
transform 1 0 14996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _530_
timestamp 1629722742
transform 1 0 14352 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_13_155
timestamp 1629722742
transform 1 0 15364 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_155
timestamp 1629722742
transform 1 0 15364 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1629722742
transform -1 0 15732 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1629722742
transform -1 0 15732 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1629722742
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1629722742
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1629722742
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _329_
timestamp 1629722742
transform 1 0 2024 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_15_17
timestamp 1629722742
transform 1 0 2668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_25
timestamp 1629722742
transform 1 0 3404 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_29
timestamp 1629722742
transform 1 0 3772 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _310_
timestamp 1629722742
transform -1 0 4784 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _311_
timestamp 1629722742
transform 1 0 3496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_40
timestamp 1629722742
transform 1 0 4784 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_46
timestamp 1629722742
transform 1 0 5336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _350_
timestamp 1629722742
transform 1 0 5428 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1629722742
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_60
timestamp 1629722742
transform 1 0 6624 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1629722742
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _309_
timestamp 1629722742
transform 1 0 6992 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _313_
timestamp 1629722742
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_71
timestamp 1629722742
transform 1 0 7636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _354_
timestamp 1629722742
transform 1 0 8004 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_81
timestamp 1629722742
transform 1 0 8556 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_87
timestamp 1629722742
transform 1 0 9108 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _274_
timestamp 1629722742
transform 1 0 9200 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1629722742
transform 1 0 9936 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _270_
timestamp 1629722742
transform -1 0 10764 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1629722742
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1629722742
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1629722742
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _478_
timestamp 1629722742
transform -1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_116
timestamp 1629722742
transform 1 0 11776 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1629722742
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _477_
timestamp 1629722742
transform -1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1629722742
transform 1 0 13248 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1629722742
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _470_
timestamp 1629722742
transform -1 0 13248 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _548_
timestamp 1629722742
transform 1 0 13616 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_148
timestamp 1629722742
transform 1 0 14720 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _285_
timestamp 1629722742
transform -1 0 14720 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1629722742
transform -1 0 15732 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_12
timestamp 1629722742
transform 1 0 2208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1629722742
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1629722742
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _331_
timestamp 1629722742
transform 1 0 1472 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1629722742
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _352_
timestamp 1629722742
transform -1 0 3220 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1629722742
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_37
timestamp 1629722742
transform 1 0 4508 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1629722742
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _314_
timestamp 1629722742
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _286_
timestamp 1629722742
transform -1 0 5888 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_16_52
timestamp 1629722742
transform 1 0 5888 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_58
timestamp 1629722742
transform 1 0 6440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _284_
timestamp 1629722742
transform 1 0 6532 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_66
timestamp 1629722742
transform 1 0 7176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _308_
timestamp 1629722742
transform 1 0 7544 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1629722742
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_88
timestamp 1629722742
transform 1 0 9200 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1629722742
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _292_
timestamp 1629722742
transform -1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_100
timestamp 1629722742
transform 1 0 10304 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_94
timestamp 1629722742
transform 1 0 9752 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _273_
timestamp 1629722742
transform 1 0 9844 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_16_106
timestamp 1629722742
transform 1 0 10856 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_113
timestamp 1629722742
transform 1 0 11500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _509_
timestamp 1629722742
transform -1 0 11500 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_122
timestamp 1629722742
transform 1 0 12328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _537_
timestamp 1629722742
transform 1 0 11868 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _550_
timestamp 1629722742
transform 1 0 12696 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1629722742
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1629722742
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1629722742
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _540_
timestamp 1629722742
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_149
timestamp 1629722742
transform 1 0 14812 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_155
timestamp 1629722742
transform 1 0 15364 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1629722742
transform -1 0 15732 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1629722742
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1629722742
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _332_
timestamp 1629722742
transform 1 0 1656 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_14
timestamp 1629722742
transform 1 0 2392 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_26
timestamp 1629722742
transform 1 0 3496 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_31
timestamp 1629722742
transform 1 0 3956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _287_
timestamp 1629722742
transform -1 0 4784 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _360_
timestamp 1629722742
transform 1 0 3588 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_40
timestamp 1629722742
transform 1 0 4784 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _330_
timestamp 1629722742
transform 1 0 5152 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1629722742
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1629722742
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1629722742
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _268_
timestamp 1629722742
transform 1 0 6716 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_67
timestamp 1629722742
transform 1 0 7268 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_76
timestamp 1629722742
transform 1 0 8096 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _482_
timestamp 1629722742
transform 1 0 7820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 1629722742
transform 1 0 8924 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _283_
timestamp 1629722742
transform 1 0 8464 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _476_
timestamp 1629722742
transform 1 0 9292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_101
timestamp 1629722742
transform 1 0 10396 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_92
timestamp 1629722742
transform 1 0 9568 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _487_
timestamp 1629722742
transform -1 0 10396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1629722742
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1629722742
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _479_
timestamp 1629722742
transform -1 0 11040 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _508_
timestamp 1629722742
transform 1 0 11500 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_17_120
timestamp 1629722742
transform 1 0 12144 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_126
timestamp 1629722742
transform 1 0 12696 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _539_
timestamp 1629722742
transform -1 0 13524 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_135
timestamp 1629722742
transform 1 0 13524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _475_
timestamp 1629722742
transform 1 0 14076 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1629722742
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_152
timestamp 1629722742
transform 1 0 15088 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1629722742
transform -1 0 15088 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1629722742
transform -1 0 15732 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1629722742
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1629722742
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1629722742
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1629722742
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_36
timestamp 1629722742
transform 1 0 4416 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1629722742
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _315_
timestamp 1629722742
transform 1 0 3772 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_44
timestamp 1629722742
transform 1 0 5152 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_1  _288_
timestamp 1629722742
transform 1 0 5336 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_54
timestamp 1629722742
transform 1 0 6072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_58
timestamp 1629722742
transform 1 0 6440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_62
timestamp 1629722742
transform 1 0 6808 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _481_
timestamp 1629722742
transform 1 0 6532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_73
timestamp 1629722742
transform 1 0 7820 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _492_
timestamp 1629722742
transform -1 0 8464 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _551_
timestamp 1629722742
transform 1 0 7176 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1629722742
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1629722742
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1629722742
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _488_
timestamp 1629722742
transform 1 0 9200 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_18_95
timestamp 1629722742
transform 1 0 9844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _489_
timestamp 1629722742
transform 1 0 10212 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_18_106
timestamp 1629722742
transform 1 0 10856 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_112
timestamp 1629722742
transform 1 0 11408 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _505_
timestamp 1629722742
transform 1 0 11500 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_18_118
timestamp 1629722742
transform 1 0 11960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_127
timestamp 1629722742
transform 1 0 12788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _538_
timestamp 1629722742
transform 1 0 12328 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1629722742
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1629722742
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1629722742
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _498_
timestamp 1629722742
transform 1 0 13156 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_18_152
timestamp 1629722742
transform 1 0 15088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _500_
timestamp 1629722742
transform -1 0 15088 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1629722742
transform -1 0 15732 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1629722742
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1629722742
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1629722742
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1629722742
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _333_
timestamp 1629722742
transform -1 0 2300 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _338_
timestamp 1629722742
transform -1 0 2760 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_19_13
timestamp 1629722742
transform 1 0 2300 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp 1629722742
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _301_
timestamp 1629722742
transform -1 0 3588 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1629722742
transform 1 0 3588 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1629722742
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1629722742
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1629722742
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _300_
timestamp 1629722742
transform 1 0 3956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_39
timestamp 1629722742
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_47
timestamp 1629722742
transform 1 0 5428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_49
timestamp 1629722742
transform 1 0 5612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_1  _303_
timestamp 1629722742
transform -1 0 5612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _517_
timestamp 1629722742
transform -1 0 5888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1629722742
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1629722742
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_62
timestamp 1629722742
transform 1 0 6808 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_61
timestamp 1629722742
transform 1 0 6716 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1629722742
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _269_
timestamp 1629722742
transform 1 0 6900 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _480_
timestamp 1629722742
transform 1 0 6532 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_68
timestamp 1629722742
transform 1 0 7360 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_69
timestamp 1629722742
transform 1 0 7452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _289_
timestamp 1629722742
transform 1 0 7820 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _519_
timestamp 1629722742
transform 1 0 7452 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_19_79
timestamp 1629722742
transform 1 0 8372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_85
timestamp 1629722742
transform 1 0 8924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1629722742
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1629722742
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _275_
timestamp 1629722742
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2b_1  _490_
timestamp 1629722742
transform -1 0 9476 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_19_91
timestamp 1629722742
transform 1 0 9476 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_95
timestamp 1629722742
transform 1 0 9844 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_93
timestamp 1629722742
transform 1 0 9660 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_99
timestamp 1629722742
transform 1 0 10212 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _493_
timestamp 1629722742
transform -1 0 10580 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _507_
timestamp 1629722742
transform -1 0 10580 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1629722742
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1629722742
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_103
timestamp 1629722742
transform 1 0 10580 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1629722742
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1629722742
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _494_
timestamp 1629722742
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _510_
timestamp 1629722742
transform -1 0 11408 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_19_119
timestamp 1629722742
transform 1 0 12052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_126
timestamp 1629722742
transform 1 0 12696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_116
timestamp 1629722742
transform 1 0 11776 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_125
timestamp 1629722742
transform 1 0 12604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _497_
timestamp 1629722742
transform 1 0 12420 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _511_
timestamp 1629722742
transform -1 0 12604 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_130
timestamp 1629722742
transform 1 0 13064 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_137
timestamp 1629722742
transform 1 0 13708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_134
timestamp 1629722742
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_141
timestamp 1629722742
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1629722742
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _495_
timestamp 1629722742
transform 1 0 13156 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _499_
timestamp 1629722742
transform -1 0 14812 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _504_
timestamp 1629722742
transform 1 0 12972 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_19_149
timestamp 1629722742
transform 1 0 14812 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_149
timestamp 1629722742
transform 1 0 14812 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _501_
timestamp 1629722742
transform -1 0 14812 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_19_155
timestamp 1629722742
transform 1 0 15364 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_155
timestamp 1629722742
transform 1 0 15364 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1629722742
transform -1 0 15732 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1629722742
transform -1 0 15732 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_11
timestamp 1629722742
transform 1 0 2116 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1629722742
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1629722742
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1629722742
transform 1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_23
timestamp 1629722742
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_1  _334_
timestamp 1629722742
transform -1 0 3220 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_35
timestamp 1629722742
transform 1 0 4324 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_39
timestamp 1629722742
transform 1 0 4692 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_48
timestamp 1629722742
transform 1 0 5520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _302_
timestamp 1629722742
transform 1 0 4784 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 1629722742
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1629722742
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _518_
timestamp 1629722742
transform 1 0 6900 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_66
timestamp 1629722742
transform 1 0 7176 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_72
timestamp 1629722742
transform 1 0 7728 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _276_
timestamp 1629722742
transform 1 0 7820 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_81
timestamp 1629722742
transform 1 0 8556 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1629722742
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1629722742
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _520_
timestamp 1629722742
transform 1 0 9476 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _546_
timestamp 1629722742
transform 1 0 10304 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1629722742
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1629722742
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1629722742
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _522_
timestamp 1629722742
transform -1 0 11776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_116
timestamp 1629722742
transform 1 0 11776 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1629722742
transform 1 0 12420 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _512_
timestamp 1629722742
transform -1 0 13524 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _525_
timestamp 1629722742
transform 1 0 12144 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_135
timestamp 1629722742
transform 1 0 13524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _483_
timestamp 1629722742
transform 1 0 14076 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_144
timestamp 1629722742
transform 1 0 14352 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_152
timestamp 1629722742
transform 1 0 15088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output25
timestamp 1629722742
transform 1 0 14720 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1629722742
transform -1 0 15732 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1629722742
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1629722742
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _365_
timestamp 1629722742
transform 1 0 1656 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_14
timestamp 1629722742
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1629722742
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_29
timestamp 1629722742
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1629722742
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _307_
timestamp 1629722742
transform 1 0 4508 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1629722742
transform 1 0 5152 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_56
timestamp 1629722742
transform 1 0 6256 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _277_
timestamp 1629722742
transform 1 0 6992 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_72
timestamp 1629722742
transform 1 0 7728 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _521_
timestamp 1629722742
transform -1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1629722742
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1629722742
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1629722742
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _549_
timestamp 1629722742
transform -1 0 9384 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_22_90
timestamp 1629722742
transform 1 0 9384 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1629722742
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _484_
timestamp 1629722742
transform -1 0 10028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _541_
timestamp 1629722742
transform 1 0 10396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_109
timestamp 1629722742
transform 1 0 11132 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_115
timestamp 1629722742
transform 1 0 11684 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1629722742
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _516_
timestamp 1629722742
transform -1 0 13064 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _526_
timestamp 1629722742
transform 1 0 11776 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_130
timestamp 1629722742
transform 1 0 13064 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1629722742
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1629722742
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _515_
timestamp 1629722742
transform 1 0 14076 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_22_148
timestamp 1629722742
transform 1 0 14720 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1629722742
transform -1 0 15732 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_10
timestamp 1629722742
transform 1 0 2024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1629722742
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _394_
timestamp 1629722742
transform 1 0 1380 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_23_18
timestamp 1629722742
transform 1 0 2760 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_24
timestamp 1629722742
transform 1 0 3312 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _335_
timestamp 1629722742
transform 1 0 3404 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output31
timestamp 1629722742
transform -1 0 2760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_33
timestamp 1629722742
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2oi_1  _305_
timestamp 1629722742
transform -1 0 5888 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1629722742
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1629722742
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1629722742
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_72
timestamp 1629722742
transform 1 0 7728 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _282_
timestamp 1629722742
transform 1 0 7084 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1629722742
transform 1 0 8832 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _280_
timestamp 1629722742
transform -1 0 9844 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_23_95
timestamp 1629722742
transform 1 0 9844 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1629722742
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1629722742
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1629722742
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1629722742
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _545_
timestamp 1629722742
transform 1 0 11592 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_121
timestamp 1629722742
transform 1 0 12236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_125
timestamp 1629722742
transform 1 0 12604 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _544_
timestamp 1629722742
transform -1 0 13340 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_133
timestamp 1629722742
transform 1 0 13340 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_137
timestamp 1629722742
transform 1 0 13708 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _513_
timestamp 1629722742
transform -1 0 14536 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_146
timestamp 1629722742
transform 1 0 14536 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_154
timestamp 1629722742
transform 1 0 15272 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1629722742
transform -1 0 15732 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_11
timestamp 1629722742
transform 1 0 2116 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1629722742
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1629722742
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _366_
timestamp 1629722742
transform 1 0 1472 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1629722742
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _336_
timestamp 1629722742
transform 1 0 2668 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1629722742
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1629722742
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _306_
timestamp 1629722742
transform 1 0 4508 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_44
timestamp 1629722742
transform 1 0 5152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _304_
timestamp 1629722742
transform 1 0 5520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1629722742
transform 1 0 6256 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_68
timestamp 1629722742
transform 1 0 7360 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1629722742
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _278_
timestamp 1629722742
transform -1 0 8188 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1629722742
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_85
timestamp 1629722742
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_89
timestamp 1629722742
transform 1 0 9292 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1629722742
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_98
timestamp 1629722742
transform 1 0 10120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _279_
timestamp 1629722742
transform 1 0 9384 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _542_
timestamp 1629722742
transform -1 0 11224 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1629722742
transform 1 0 11224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1629722742
transform 1 0 11592 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_117
timestamp 1629722742
transform 1 0 11868 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _543_
timestamp 1629722742
transform -1 0 12972 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_129
timestamp 1629722742
transform 1 0 12972 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1629722742
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_141
timestamp 1629722742
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1629722742
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _531_
timestamp 1629722742
transform -1 0 13616 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_151
timestamp 1629722742
transform 1 0 14996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _514_
timestamp 1629722742
transform -1 0 14996 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_24_155
timestamp 1629722742
transform 1 0 15364 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1629722742
transform -1 0 15732 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1629722742
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1629722742
transform 1 0 1380 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_25_13
timestamp 1629722742
transform 1 0 2300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_24
timestamp 1629722742
transform 1 0 3312 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _337_
timestamp 1629722742
transform 1 0 2668 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_25_29
timestamp 1629722742
transform 1 0 3772 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_37
timestamp 1629722742
transform 1 0 4508 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1629722742
transform 1 0 3680 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output18
timestamp 1629722742
transform -1 0 4508 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1629722742
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output22
timestamp 1629722742
transform -1 0 5244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1629722742
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1629722742
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1629722742
transform 1 0 6348 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_25_67
timestamp 1629722742
transform 1 0 7268 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_75
timestamp 1629722742
transform 1 0 8004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output27
timestamp 1629722742
transform -1 0 8004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_83
timestamp 1629722742
transform 1 0 8740 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1629722742
transform 1 0 8832 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _281_
timestamp 1629722742
transform 1 0 8924 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_25_100
timestamp 1629722742
transform 1 0 10304 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_92
timestamp 1629722742
transform 1 0 9568 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output28
timestamp 1629722742
transform -1 0 10304 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1629722742
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1629722742
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_116
timestamp 1629722742
transform 1 0 11776 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_127
timestamp 1629722742
transform 1 0 12788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1629722742
transform -1 0 12788 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1629722742
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_139
timestamp 1629722742
transform 1 0 13892 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1629722742
transform 1 0 13984 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _533_
timestamp 1629722742
transform -1 0 14352 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1629722742
transform 1 0 13156 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_144
timestamp 1629722742
transform 1 0 14352 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1629722742
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output26
timestamp 1629722742
transform 1 0 14720 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1629722742
transform -1 0 15732 0 -1 16320
box -38 -48 314 592
<< labels >>
rlabel metal5 s 1104 6682 15732 7002 4 VGND
port 1 nsew
rlabel metal5 s 1104 4326 15732 4646 4 VPWR
port 2 nsew
rlabel metal2 s 16762 18215 16818 19015 4 a[0]
port 3 nsew
rlabel metal3 s 0 16328 800 16448 4 a[1]
port 4 nsew
rlabel metal3 s 0 5448 800 5568 4 a[2]
port 5 nsew
rlabel metal2 s 7378 0 7434 800 4 a[3]
port 6 nsew
rlabel metal2 s 5722 18215 5778 19015 4 a[4]
port 7 nsew
rlabel metal2 s 11242 18215 11298 19015 4 a[5]
port 8 nsew
rlabel metal2 s 12898 0 12954 800 4 a[6]
port 9 nsew
rlabel metal3 s 16071 7896 16871 8016 4 a[7]
port 10 nsew
rlabel metal2 s 11058 0 11114 800 4 b[0]
port 11 nsew
rlabel metal3 s 16071 10616 16871 10736 4 b[1]
port 12 nsew
rlabel metal3 s 0 2728 800 2848 4 b[2]
port 13 nsew
rlabel metal2 s 18 0 74 800 4 b[3]
port 14 nsew
rlabel metal2 s 13082 18215 13138 19015 4 b[4]
port 15 nsew
rlabel metal2 s 14922 18215 14978 19015 4 b[5]
port 16 nsew
rlabel metal3 s 0 13608 800 13728 4 b[6]
port 17 nsew
rlabel metal2 s 16762 0 16818 800 4 b[7]
port 18 nsew
rlabel metal3 s 0 8168 800 8288 4 m[0]
port 19 nsew
rlabel metal2 s 18 18215 74 19015 4 m[10]
port 20 nsew
rlabel metal2 s 14922 0 14978 800 4 m[11]
port 21 nsew
rlabel metal2 s 1858 0 1914 800 4 m[12]
port 22 nsew
rlabel metal2 s 3698 0 3754 800 4 m[13]
port 23 nsew
rlabel metal2 s 3882 18215 3938 19015 4 m[14]
port 24 nsew
rlabel metal3 s 16071 2456 16871 2576 4 m[15]
port 25 nsew
rlabel metal2 s 5538 0 5594 800 4 m[1]
port 26 nsew
rlabel metal3 s 16071 13336 16871 13456 4 m[2]
port 27 nsew
rlabel metal3 s 16071 16056 16871 16176 4 m[3]
port 28 nsew
rlabel metal2 s 7562 18215 7618 19015 4 m[4]
port 29 nsew
rlabel metal2 s 9402 18215 9458 19015 4 m[5]
port 30 nsew
rlabel metal2 s 9218 0 9274 800 4 m[6]
port 31 nsew
rlabel metal3 s 0 10888 800 11008 4 m[7]
port 32 nsew
rlabel metal2 s 1858 18215 1914 19015 4 m[8]
port 33 nsew
rlabel metal3 s 16071 5176 16871 5296 4 m[9]
port 34 nsew
<< properties >>
string FIXED_BBOX 0 0 16871 19015
<< end >>

* NGSPICE file created from dvsd_8216m9.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

.subckt dvsd_8216m9 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] B[0] B[1] B[2] B[3] B[4]
+ B[5] B[6] B[7] M[0] M[10] M[11] M[12] M[13] M[14] M[15] M[1] M[2] M[3] M[4] M[5]
+ M[6] M[7] M[8] M[9] VGND VPWR
X_432_ _432_/A _432_/B VGND VGND VPWR VPWR _432_/X sky130_fd_sc_hd__or2_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_501_ _531_/A _531_/C _531_/A _531_/C VGND VGND VPWR VPWR _501_/Y sky130_fd_sc_hd__a2bb2oi_1
X_363_ _363_/A _363_/B VGND VGND VPWR VPWR _430_/A sky130_fd_sc_hd__or2_1
XFILLER_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_346_ _346_/A VGND VGND VPWR VPWR _347_/A sky130_fd_sc_hd__buf_6
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_415_ _448_/A VGND VGND VPWR VPWR _561_/A sky130_fd_sc_hd__buf_1
X_329_ _314_/X _328_/X _314_/X _328_/X VGND VGND VPWR VPWR _329_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_594_ _573_/A _593_/Y _573_/Y _593_/A VGND VGND VPWR VPWR _594_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput31 _501_/Y VGND VGND VPWR VPWR M[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput20 _607_/X VGND VGND VPWR VPWR M[12] sky130_fd_sc_hd__clkbuf_2
X_577_ _559_/X _576_/X _559_/X _576_/X VGND VGND VPWR VPWR _580_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_431_ _428_/X _430_/X _428_/X _430_/X VGND VGND VPWR VPWR _431_/X sky130_fd_sc_hd__a2bb2o_1
X_362_ _351_/X _361_/X _351_/X _361_/X VGND VGND VPWR VPWR _363_/B sky130_fd_sc_hd__a2bb2o_1
X_500_ _427_/A _464_/A _465_/X _466_/X VGND VGND VPWR VPWR _531_/C sky130_fd_sc_hd__o22a_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_629_ _629_/A _629_/B VGND VGND VPWR VPWR _629_/X sky130_fd_sc_hd__or2_1
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_345_ _442_/B VGND VGND VPWR VPWR _346_/A sky130_fd_sc_hd__inv_2
X_414_ _542_/A VGND VGND VPWR VPWR _448_/A sky130_fd_sc_hd__inv_2
X_328_ _328_/A _328_/B VGND VGND VPWR VPWR _328_/X sky130_fd_sc_hd__or2_1
XFILLER_9_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_593_ _593_/A VGND VGND VPWR VPWR _593_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput21 _620_/X VGND VGND VPWR VPWR M[13] sky130_fd_sc_hd__clkbuf_2
X_576_ _574_/X _575_/X _574_/X _575_/X VGND VGND VPWR VPWR _576_/X sky130_fd_sc_hd__a2bb2o_1
Xoutput32 _530_/X VGND VGND VPWR VPWR M[9] sky130_fd_sc_hd__clkbuf_2
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_361_ _352_/X _360_/X _352_/X _360_/X VGND VGND VPWR VPWR _361_/X sky130_fd_sc_hd__a2bb2o_1
X_430_ _430_/A _432_/B VGND VGND VPWR VPWR _430_/X sky130_fd_sc_hd__or2_1
XFILLER_13_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_628_ _621_/X _622_/X _623_/X _625_/Y _627_/X VGND VGND VPWR VPWR _628_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_559_ _570_/A _503_/A _535_/Y _538_/Y _539_/X VGND VGND VPWR VPWR _559_/X sky130_fd_sc_hd__o32a_1
XFILLER_12_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_344_ _329_/X _338_/X _342_/X _343_/X VGND VGND VPWR VPWR _363_/A sky130_fd_sc_hd__o22a_1
X_413_ _447_/B _516_/A VGND VGND VPWR VPWR _413_/X sky130_fd_sc_hd__or2_1
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_327_ _631_/A _481_/A _367_/C _445_/A VGND VGND VPWR VPWR _328_/B sky130_fd_sc_hd__o22a_1
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_592_ _590_/A _590_/B _591_/Y VGND VGND VPWR VPWR _593_/A sky130_fd_sc_hd__a21oi_1
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput22 _626_/Y VGND VGND VPWR VPWR M[14] sky130_fd_sc_hd__clkbuf_2
X_575_ _546_/X _547_/X _540_/X _548_/X VGND VGND VPWR VPWR _575_/X sky130_fd_sc_hd__o22a_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ _353_/X _359_/X _353_/X _359_/X VGND VGND VPWR VPWR _360_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_558_ _557_/A _557_/B _556_/Y _556_/A _557_/Y VGND VGND VPWR VPWR _558_/X sky130_fd_sc_hd__o32a_1
X_489_ _483_/X _488_/X _483_/X _488_/X VGND VGND VPWR VPWR _489_/X sky130_fd_sc_hd__a2bb2o_1
X_627_ _627_/A _627_/B _627_/C _627_/D VGND VGND VPWR VPWR _627_/X sky130_fd_sc_hd__or4_1
XFILLER_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_343_ _329_/X _338_/X _329_/X _338_/X VGND VGND VPWR VPWR _343_/X sky130_fd_sc_hd__a2bb2o_1
X_412_ _408_/X _411_/X _408_/X _411_/X VGND VGND VPWR VPWR _412_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_326_ _326_/A VGND VGND VPWR VPWR _445_/A sky130_fd_sc_hd__buf_1
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_591_ _591_/A VGND VGND VPWR VPWR _591_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput23 _628_/Y VGND VGND VPWR VPWR M[15] sky130_fd_sc_hd__clkbuf_2
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_574_ _572_/A _572_/B _573_/Y VGND VGND VPWR VPWR _574_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_557_ _557_/A _557_/B VGND VGND VPWR VPWR _557_/Y sky130_fd_sc_hd__nor2_1
X_626_ _623_/X _625_/Y _623_/X _625_/Y VGND VGND VPWR VPWR _626_/Y sky130_fd_sc_hd__a2bb2oi_1
X_488_ _486_/X _487_/X _486_/X _487_/X VGND VGND VPWR VPWR _488_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_342_ _350_/C _631_/B VGND VGND VPWR VPWR _342_/X sky130_fd_sc_hd__or2_1
X_411_ _411_/A _411_/B VGND VGND VPWR VPWR _411_/X sky130_fd_sc_hd__or2_1
XFILLER_12_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_609_ _542_/D _469_/X _622_/C _608_/X VGND VGND VPWR VPWR _610_/A sky130_fd_sc_hd__a31o_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_325_ _390_/D VGND VGND VPWR VPWR _326_/A sky130_fd_sc_hd__inv_2
XFILLER_18_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_590_ _590_/A _590_/B VGND VGND VPWR VPWR _591_/A sky130_fd_sc_hd__or2_1
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput24 _633_/Y VGND VGND VPWR VPWR M[1] sky130_fd_sc_hd__clkbuf_2
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_573_ _573_/A VGND VGND VPWR VPWR _573_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_625_ _601_/A _618_/A _606_/A _624_/X VGND VGND VPWR VPWR _625_/Y sky130_fd_sc_hd__a31oi_2
X_556_ _556_/A VGND VGND VPWR VPWR _556_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_487_ _449_/A _452_/X _447_/X _453_/X VGND VGND VPWR VPWR _487_/X sky130_fd_sc_hd__o22a_1
X_341_ _436_/A VGND VGND VPWR VPWR _631_/B sky130_fd_sc_hd__buf_1
X_410_ _542_/B _410_/B _410_/C _542_/C VGND VGND VPWR VPWR _411_/B sky130_fd_sc_hd__and4_1
XFILLER_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_539_ _539_/A _587_/A VGND VGND VPWR VPWR _539_/X sky130_fd_sc_hd__or2_1
X_608_ _627_/A _627_/B _627_/C _627_/D VGND VGND VPWR VPWR _608_/X sky130_fd_sc_hd__o22a_1
XFILLER_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_324_ _448_/B VGND VGND VPWR VPWR _367_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput25 _634_/Y VGND VGND VPWR VPWR M[2] sky130_fd_sc_hd__clkbuf_2
X_572_ _572_/A _572_/B VGND VGND VPWR VPWR _573_/A sky130_fd_sc_hd__or2_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_555_ _554_/A _554_/B _554_/X VGND VGND VPWR VPWR _556_/A sky130_fd_sc_hd__a21bo_1
X_624_ _616_/A _616_/B _599_/Y _616_/Y VGND VGND VPWR VPWR _624_/X sky130_fd_sc_hd__o2bb2a_1
X_486_ _486_/A _486_/B VGND VGND VPWR VPWR _486_/X sky130_fd_sc_hd__or2_1
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_340_ _340_/A VGND VGND VPWR VPWR _350_/C sky130_fd_sc_hd__clkbuf_2
X_607_ _601_/Y _606_/Y _601_/A _606_/A VGND VGND VPWR VPWR _607_/X sky130_fd_sc_hd__o22a_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_538_ _538_/A VGND VGND VPWR VPWR _538_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_469_ _469_/A VGND VGND VPWR VPWR _469_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_323_ _417_/A VGND VGND VPWR VPWR _448_/B sky130_fd_sc_hd__inv_2
XFILLER_1_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput26 _635_/Y VGND VGND VPWR VPWR M[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_571_ _381_/B _469_/X _569_/A _569_/Y _570_/X VGND VGND VPWR VPWR _572_/B sky130_fd_sc_hd__a32o_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_554_ _554_/A _554_/B VGND VGND VPWR VPWR _554_/X sky130_fd_sc_hd__or2_1
X_623_ _621_/X _622_/X _621_/X _622_/X VGND VGND VPWR VPWR _623_/X sky130_fd_sc_hd__a2bb2o_1
X_485_ _485_/A _542_/D _542_/A _485_/D VGND VGND VPWR VPWR _486_/B sky130_fd_sc_hd__and4_1
X_399_ _374_/X _397_/X _350_/X _398_/X VGND VGND VPWR VPWR _426_/A sky130_fd_sc_hd__o22a_1
XFILLER_27_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_468_ _437_/X _438_/X _436_/X _439_/X VGND VGND VPWR VPWR _468_/X sky130_fd_sc_hd__o22a_1
XFILLER_4_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_606_ _606_/A VGND VGND VPWR VPWR _606_/Y sky130_fd_sc_hd__inv_2
X_537_ _570_/A _472_/B _535_/Y _535_/A _536_/Y VGND VGND VPWR VPWR _538_/A sky130_fd_sc_hd__o32a_1
XFILLER_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_322_ _322_/A VGND VGND VPWR VPWR _481_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput27 _373_/Y VGND VGND VPWR VPWR M[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_570_ _570_/A _570_/B VGND VGND VPWR VPWR _570_/X sky130_fd_sc_hd__or2_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_553_ _523_/X _524_/X _504_/X _525_/X VGND VGND VPWR VPWR _554_/B sky130_fd_sc_hd__o22a_1
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_622_ _627_/B _627_/D _622_/C VGND VGND VPWR VPWR _622_/X sky130_fd_sc_hd__or3_1
X_484_ _367_/C _563_/B _561_/A _519_/A VGND VGND VPWR VPWR _486_/A sky130_fd_sc_hd__o22a_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_398_ _374_/X _397_/X _374_/X _397_/X VGND VGND VPWR VPWR _398_/X sky130_fd_sc_hd__a2bb2o_1
X_467_ _465_/X _466_/X _465_/X _466_/X VGND VGND VPWR VPWR _467_/Y sky130_fd_sc_hd__a2bb2oi_1
X_605_ _556_/Y _602_/Y _557_/A _604_/X VGND VGND VPWR VPWR _606_/A sky130_fd_sc_hd__a31o_1
X_536_ _570_/A _585_/B VGND VGND VPWR VPWR _536_/Y sky130_fd_sc_hd__nor2_1
X_321_ _442_/A VGND VGND VPWR VPWR _322_/A sky130_fd_sc_hd__inv_2
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_519_ _519_/A _563_/B _519_/C VGND VGND VPWR VPWR _519_/X sky130_fd_sc_hd__or3_1
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput28 _630_/X VGND VGND VPWR VPWR M[5] sky130_fd_sc_hd__clkbuf_2
Xoutput17 _631_/Y VGND VGND VPWR VPWR M[0] sky130_fd_sc_hd__clkbuf_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_552_ _533_/X _551_/X _533_/X _551_/X VGND VGND VPWR VPWR _554_/A sky130_fd_sc_hd__a2bb2o_1
X_483_ _410_/C _386_/X _480_/Y _482_/X _480_/A VGND VGND VPWR VPWR _483_/X sky130_fd_sc_hd__a32o_1
X_621_ _591_/A _610_/A _611_/X _613_/X VGND VGND VPWR VPWR _621_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_466_ _428_/X _430_/X _431_/X _432_/X VGND VGND VPWR VPWR _466_/X sky130_fd_sc_hd__o22a_1
X_397_ _384_/X _396_/X _384_/X _396_/X VGND VGND VPWR VPWR _397_/X sky130_fd_sc_hd__a2bb2o_1
X_604_ _556_/Y _602_/Y _557_/B _603_/Y VGND VGND VPWR VPWR _604_/X sky130_fd_sc_hd__a31o_1
X_535_ _535_/A VGND VGND VPWR VPWR _535_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_320_ _452_/A VGND VGND VPWR VPWR _631_/A sky130_fd_sc_hd__buf_6
XFILLER_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_449_ _449_/A VGND VGND VPWR VPWR _519_/C sky130_fd_sc_hd__inv_2
X_518_ _381_/B _386_/X _515_/Y _517_/X _515_/A VGND VGND VPWR VPWR _518_/X sky130_fd_sc_hd__a32o_1
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput18 _558_/X VGND VGND VPWR VPWR M[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput29 _433_/Y VGND VGND VPWR VPWR M[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_24_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_620_ _618_/Y _619_/Y _618_/Y _619_/Y VGND VGND VPWR VPWR _620_/X sky130_fd_sc_hd__a2bb2o_1
X_551_ _549_/X _550_/X _549_/X _550_/X VGND VGND VPWR VPWR _551_/X sky130_fd_sc_hd__a2bb2o_1
X_482_ _539_/A _563_/D VGND VGND VPWR VPWR _482_/X sky130_fd_sc_hd__or2_1
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_465_ _427_/A _464_/A _427_/Y _464_/Y VGND VGND VPWR VPWR _465_/X sky130_fd_sc_hd__a22o_1
X_396_ _386_/X _330_/A _392_/Y _395_/X _392_/A VGND VGND VPWR VPWR _396_/X sky130_fd_sc_hd__a32o_1
X_603_ _554_/X _579_/X _581_/B VGND VGND VPWR VPWR _603_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_534_ _381_/B _386_/A _515_/Y _514_/B VGND VGND VPWR VPWR _535_/A sky130_fd_sc_hd__a31o_1
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_448_ _448_/A _448_/B VGND VGND VPWR VPWR _449_/A sky130_fd_sc_hd__or2_1
X_517_ _570_/A _584_/A VGND VGND VPWR VPWR _517_/X sky130_fd_sc_hd__or2_1
X_379_ _448_/B _516_/A _452_/A _544_/A VGND VGND VPWR VPWR _382_/A sky130_fd_sc_hd__o22a_1
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput19 _583_/X VGND VGND VPWR VPWR M[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_481_ _481_/A VGND VGND VPWR VPWR _539_/A sky130_fd_sc_hd__buf_1
X_550_ _520_/X _521_/X _511_/X _522_/X VGND VGND VPWR VPWR _550_/X sky130_fd_sc_hd__o22a_1
XFILLER_27_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_464_ _464_/A VGND VGND VPWR VPWR _464_/Y sky130_fd_sc_hd__inv_2
X_602_ _602_/A VGND VGND VPWR VPWR _602_/Y sky130_fd_sc_hd__inv_2
X_533_ _539_/A _503_/A _506_/Y _509_/Y _510_/X VGND VGND VPWR VPWR _533_/X sky130_fd_sc_hd__o32a_1
X_395_ _584_/A _436_/A VGND VGND VPWR VPWR _395_/X sky130_fd_sc_hd__or2_1
X_378_ _378_/A VGND VGND VPWR VPWR _544_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_447_ _544_/A _447_/B VGND VGND VPWR VPWR _447_/X sky130_fd_sc_hd__or2_1
X_516_ _516_/A VGND VGND VPWR VPWR _570_/A sky130_fd_sc_hd__buf_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_480_ _480_/A VGND VGND VPWR VPWR _480_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_601_ _601_/A VGND VGND VPWR VPWR _601_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_463_ _406_/Y _462_/X _406_/Y _462_/X VGND VGND VPWR VPWR _464_/A sky130_fd_sc_hd__a2bb2o_1
X_532_ _527_/A _527_/B _498_/Y _527_/Y VGND VGND VPWR VPWR _557_/B sky130_fd_sc_hd__o2bb2a_1
X_394_ _563_/D VGND VGND VPWR VPWR _584_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_446_ _410_/B _386_/X _444_/Y _445_/X _444_/A VGND VGND VPWR VPWR _446_/X sky130_fd_sc_hd__a32o_1
XFILLER_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_377_ _380_/A VGND VGND VPWR VPWR _378_/A sky130_fd_sc_hd__inv_2
X_515_ _515_/A VGND VGND VPWR VPWR _515_/Y sky130_fd_sc_hd__inv_2
X_429_ _350_/X _398_/X _350_/X _398_/X VGND VGND VPWR VPWR _432_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 A[0] VGND VGND VPWR VPWR _330_/A sky130_fd_sc_hd__buf_1
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_531_ _531_/A _531_/B _531_/C VGND VGND VPWR VPWR _557_/A sky130_fd_sc_hd__nor3_1
X_462_ _460_/X _461_/X _460_/X _461_/X VGND VGND VPWR VPWR _462_/X sky130_fd_sc_hd__a2bb2o_1
X_393_ _393_/A VGND VGND VPWR VPWR _563_/D sky130_fd_sc_hd__inv_2
XFILLER_4_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_600_ _598_/A _598_/B _599_/Y VGND VGND VPWR VPWR _601_/A sky130_fd_sc_hd__a21oi_2
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_514_ _514_/A _514_/B VGND VGND VPWR VPWR _515_/A sky130_fd_sc_hd__or2_1
X_445_ _445_/A _563_/D VGND VGND VPWR VPWR _445_/X sky130_fd_sc_hd__or2_1
X_376_ _447_/B _481_/A VGND VGND VPWR VPWR _376_/X sky130_fd_sc_hd__or2_1
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_428_ _426_/A _426_/B _427_/Y VGND VGND VPWR VPWR _428_/X sky130_fd_sc_hd__a21o_1
X_359_ _359_/A _359_/B VGND VGND VPWR VPWR _359_/X sky130_fd_sc_hd__or2_1
Xinput2 A[1] VGND VGND VPWR VPWR _390_/B sky130_fd_sc_hd__clkbuf_2
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_530_ _531_/B _529_/Y _531_/B _529_/Y VGND VGND VPWR VPWR _530_/X sky130_fd_sc_hd__a2bb2o_1
X_461_ _422_/X _423_/X _407_/Y _424_/X VGND VGND VPWR VPWR _461_/X sky130_fd_sc_hd__o22a_1
X_392_ _392_/A VGND VGND VPWR VPWR _392_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_444_ _444_/A VGND VGND VPWR VPWR _444_/Y sky130_fd_sc_hd__inv_2
X_375_ _353_/X _359_/X _359_/B VGND VGND VPWR VPWR _375_/X sky130_fd_sc_hd__o21ba_1
X_513_ _513_/A _542_/B _542_/A _542_/C VGND VGND VPWR VPWR _514_/B sky130_fd_sc_hd__and4_1
X_427_ _427_/A VGND VGND VPWR VPWR _427_/Y sky130_fd_sc_hd__inv_2
X_358_ _485_/A _442_/A _381_/C _381_/B VGND VGND VPWR VPWR _359_/B sky130_fd_sc_hd__and4_1
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 A[2] VGND VGND VPWR VPWR _390_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_391_ _391_/A _391_/B VGND VGND VPWR VPWR _392_/A sky130_fd_sc_hd__or2_1
X_460_ _440_/X _459_/X _440_/X _459_/X VGND VGND VPWR VPWR _460_/X sky130_fd_sc_hd__a2bb2o_1
X_589_ _612_/A _588_/Y _612_/A _588_/Y VGND VGND VPWR VPWR _590_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_374_ _352_/X _360_/X _351_/X _361_/X VGND VGND VPWR VPWR _374_/X sky130_fd_sc_hd__o22a_1
X_443_ _443_/A _443_/B VGND VGND VPWR VPWR _444_/A sky130_fd_sc_hd__or2_1
X_512_ _378_/A _347_/A _561_/A _340_/A VGND VGND VPWR VPWR _514_/A sky130_fd_sc_hd__o22a_1
XFILLER_24_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_426_ _426_/A _426_/B VGND VGND VPWR VPWR _427_/A sky130_fd_sc_hd__or2_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_357_ _478_/A VGND VGND VPWR VPWR _381_/B sky130_fd_sc_hd__clkbuf_2
Xinput4 A[3] VGND VGND VPWR VPWR _442_/A sky130_fd_sc_hd__buf_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_409_ _563_/A _326_/A _481_/A _350_/C VGND VGND VPWR VPWR _411_/A sky130_fd_sc_hd__o22a_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_390_ _542_/B _390_/B _542_/C _390_/D VGND VGND VPWR VPWR _391_/B sky130_fd_sc_hd__and4_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_588_ _588_/A _627_/D VGND VGND VPWR VPWR _588_/Y sky130_fd_sc_hd__nor2_1
X_373_ _371_/A _371_/B _629_/B VGND VGND VPWR VPWR _373_/Y sky130_fd_sc_hd__a21oi_1
X_442_ _442_/A _442_/B _478_/A _442_/D VGND VGND VPWR VPWR _443_/B sky130_fd_sc_hd__and4_1
X_511_ _410_/B _469_/X _509_/A _509_/Y _510_/X VGND VGND VPWR VPWR _511_/X sky130_fd_sc_hd__a32o_1
XFILLER_5_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput5 A[4] VGND VGND VPWR VPWR _478_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_425_ _407_/Y _424_/X _407_/Y _424_/X VGND VGND VPWR VPWR _426_/B sky130_fd_sc_hd__a2bb2o_1
X_356_ _448_/B _481_/A _452_/A _516_/A VGND VGND VPWR VPWR _359_/A sky130_fd_sc_hd__o22a_1
XFILLER_27_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ _563_/D _408_/B VGND VGND VPWR VPWR _408_/X sky130_fd_sc_hd__or2_1
X_339_ _442_/D VGND VGND VPWR VPWR _340_/A sky130_fd_sc_hd__inv_2
XFILLER_7_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_587_ _587_/A VGND VGND VPWR VPWR _627_/D sky130_fd_sc_hd__buf_1
X_372_ _432_/A VGND VGND VPWR VPWR _629_/B sky130_fd_sc_hd__inv_2
X_510_ _510_/A _587_/A VGND VGND VPWR VPWR _510_/X sky130_fd_sc_hd__or2_1
X_441_ _322_/A _346_/A _355_/A _340_/A VGND VGND VPWR VPWR _443_/A sky130_fd_sc_hd__o22a_1
XFILLER_1_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_424_ _422_/X _423_/X _422_/X _423_/X VGND VGND VPWR VPWR _424_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_355_ _355_/A VGND VGND VPWR VPWR _516_/A sky130_fd_sc_hd__buf_6
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput6 A[5] VGND VGND VPWR VPWR _380_/A sky130_fd_sc_hd__buf_1
XFILLER_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_407_ _406_/A _406_/B _406_/Y VGND VGND VPWR VPWR _407_/Y sky130_fd_sc_hd__o21ai_1
X_338_ _332_/X _337_/X _337_/A VGND VGND VPWR VPWR _338_/X sky130_fd_sc_hd__o21ba_1
XFILLER_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_586_ _503_/A _622_/C _586_/S VGND VGND VPWR VPWR _612_/A sky130_fd_sc_hd__mux2_1
X_371_ _371_/A _371_/B VGND VGND VPWR VPWR _432_/A sky130_fd_sc_hd__or2_1
X_440_ _436_/X _439_/X _436_/X _439_/X VGND VGND VPWR VPWR _440_/X sky130_fd_sc_hd__a2bb2o_1
X_569_ _569_/A VGND VGND VPWR VPWR _569_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_423_ _375_/X _383_/X _384_/X _396_/X VGND VGND VPWR VPWR _423_/X sky130_fd_sc_hd__o22a_1
X_354_ _478_/A VGND VGND VPWR VPWR _355_/A sky130_fd_sc_hd__inv_2
XFILLER_6_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 A[6] VGND VGND VPWR VPWR _542_/A sky130_fd_sc_hd__buf_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_406_ _406_/A _406_/B VGND VGND VPWR VPWR _406_/Y sky130_fd_sc_hd__nand2_1
X_337_ _337_/A _337_/B VGND VGND VPWR VPWR _337_/X sky130_fd_sc_hd__or2_1
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput10 B[1] VGND VGND VPWR VPWR _417_/A sky130_fd_sc_hd__buf_1
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_585_ _627_/C _585_/B VGND VGND VPWR VPWR _622_/C sky130_fd_sc_hd__nor2_1
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_370_ _370_/A _370_/B VGND VGND VPWR VPWR _371_/B sky130_fd_sc_hd__or2_1
X_499_ _497_/A _497_/B _498_/Y VGND VGND VPWR VPWR _531_/A sky130_fd_sc_hd__a21o_1
X_568_ _544_/A _567_/B _566_/Y _566_/A _567_/Y VGND VGND VPWR VPWR _569_/A sky130_fd_sc_hd__o32a_1
X_422_ _412_/X _421_/X _412_/X _421_/X VGND VGND VPWR VPWR _422_/X sky130_fd_sc_hd__a2bb2o_1
X_353_ _519_/A _445_/A VGND VGND VPWR VPWR _353_/X sky130_fd_sc_hd__or2_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 A[7] VGND VGND VPWR VPWR _542_/D sky130_fd_sc_hd__clkbuf_2
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_405_ _631_/B _503_/A VGND VGND VPWR VPWR _406_/B sky130_fd_sc_hd__nor2_1
X_336_ _631_/A _510_/A _367_/C _408_/B VGND VGND VPWR VPWR _337_/B sky130_fd_sc_hd__o22a_1
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_319_ _417_/D VGND VGND VPWR VPWR _452_/A sky130_fd_sc_hd__inv_2
Xinput11 B[2] VGND VGND VPWR VPWR _485_/D sky130_fd_sc_hd__buf_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_584_ _584_/A _627_/B VGND VGND VPWR VPWR _590_/A sky130_fd_sc_hd__or2_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_498_ _498_/A VGND VGND VPWR VPWR _498_/Y sky130_fd_sc_hd__inv_2
X_567_ _588_/A _567_/B VGND VGND VPWR VPWR _567_/Y sky130_fd_sc_hd__nor2_1
X_421_ _419_/X _420_/X _419_/X _420_/X VGND VGND VPWR VPWR _421_/X sky130_fd_sc_hd__a2bb2o_1
X_352_ _314_/X _328_/X _328_/A VGND VGND VPWR VPWR _352_/X sky130_fd_sc_hd__o21ba_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_619_ _601_/Y _606_/Y _599_/A VGND VGND VPWR VPWR _619_/Y sky130_fd_sc_hd__o21ai_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 B[0] VGND VGND VPWR VPWR _417_/D sky130_fd_sc_hd__buf_1
XFILLER_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_335_ _445_/A VGND VGND VPWR VPWR _510_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_404_ _585_/B VGND VGND VPWR VPWR _503_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_318_ _381_/C _410_/C _485_/A _390_/D VGND VGND VPWR VPWR _328_/A sky130_fd_sc_hd__and4_1
Xinput12 B[3] VGND VGND VPWR VPWR _442_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_583_ _602_/A _582_/Y _602_/A _582_/Y VGND VGND VPWR VPWR _583_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_635_ _370_/A _370_/B _371_/B VGND VGND VPWR VPWR _635_/Y sky130_fd_sc_hd__a21boi_1
X_497_ _497_/A _497_/B VGND VGND VPWR VPWR _498_/A sky130_fd_sc_hd__or2_1
XFILLER_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_566_ _566_/A VGND VGND VPWR VPWR _566_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_351_ _351_/A _350_/X VGND VGND VPWR VPWR _351_/X sky130_fd_sc_hd__or2b_1
X_420_ _376_/X _382_/X _382_/B VGND VGND VPWR VPWR _420_/X sky130_fd_sc_hd__o21ba_1
XFILLER_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_618_ _618_/A VGND VGND VPWR VPWR _618_/Y sky130_fd_sc_hd__inv_2
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_549_ _540_/X _548_/X _540_/X _548_/X VGND VGND VPWR VPWR _549_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_334_ _381_/C _410_/B _485_/A _390_/B VGND VGND VPWR VPWR _337_/A sky130_fd_sc_hd__and4_1
X_403_ _472_/B VGND VGND VPWR VPWR _585_/B sky130_fd_sc_hd__buf_1
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 B[4] VGND VGND VPWR VPWR _442_/B sky130_fd_sc_hd__buf_1
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_317_ _417_/A VGND VGND VPWR VPWR _485_/A sky130_fd_sc_hd__buf_1
XFILLER_20_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_582_ _556_/A _557_/Y _554_/X VGND VGND VPWR VPWR _582_/Y sky130_fd_sc_hd__o21ai_1
X_496_ _460_/X _461_/X _406_/Y _462_/X VGND VGND VPWR VPWR _497_/B sky130_fd_sc_hd__o22a_1
X_634_ _368_/A _368_/B _370_/A VGND VGND VPWR VPWR _634_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_565_ _513_/A _386_/A _543_/Y _543_/B VGND VGND VPWR VPWR _566_/A sky130_fd_sc_hd__a31o_1
XFILLER_5_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_350_ _563_/A _350_/B _350_/C _408_/B VGND VGND VPWR VPWR _350_/X sky130_fd_sc_hd__or4_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_617_ _616_/A _616_/B _616_/Y VGND VGND VPWR VPWR _618_/A sky130_fd_sc_hd__a21oi_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_548_ _546_/X _547_/X _546_/X _547_/X VGND VGND VPWR VPWR _548_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_479_ _479_/A _479_/B VGND VGND VPWR VPWR _480_/A sky130_fd_sc_hd__or2_1
XFILLER_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_402_ _567_/B VGND VGND VPWR VPWR _472_/B sky130_fd_sc_hd__buf_1
X_333_ _390_/D VGND VGND VPWR VPWR _410_/B sky130_fd_sc_hd__buf_1
Xinput14 B[5] VGND VGND VPWR VPWR _393_/A sky130_fd_sc_hd__buf_1
X_316_ _442_/A VGND VGND VPWR VPWR _410_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_581_ _579_/X _581_/B VGND VGND VPWR VPWR _602_/A sky130_fd_sc_hd__nand2b_1
XFILLER_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_495_ _468_/X _494_/X _468_/X _494_/X VGND VGND VPWR VPWR _497_/A sky130_fd_sc_hd__a2bb2o_1
X_633_ _633_/A _368_/B VGND VGND VPWR VPWR _633_/Y sky130_fd_sc_hd__nor2b_1
X_564_ _564_/A _586_/S VGND VGND VPWR VPWR _572_/A sky130_fd_sc_hd__or2b_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_478_ _478_/A _542_/B _513_/A _542_/C VGND VGND VPWR VPWR _479_/B sky130_fd_sc_hd__and4_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_616_ _616_/A _616_/B VGND VGND VPWR VPWR _616_/Y sky130_fd_sc_hd__nor2_1
X_547_ _518_/X _519_/X _486_/B VGND VGND VPWR VPWR _547_/X sky130_fd_sc_hd__o21ba_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_401_ _401_/A VGND VGND VPWR VPWR _567_/B sky130_fd_sc_hd__inv_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_332_ _519_/A _436_/A VGND VGND VPWR VPWR _332_/X sky130_fd_sc_hd__or2_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput15 B[6] VGND VGND VPWR VPWR _401_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_315_ _417_/D VGND VGND VPWR VPWR _381_/C sky130_fd_sc_hd__buf_6
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_580_ _580_/A _580_/B VGND VGND VPWR VPWR _581_/B sky130_fd_sc_hd__or2_1
X_632_ _631_/A _475_/A _367_/C _631_/B VGND VGND VPWR VPWR _633_/A sky130_fd_sc_hd__o22a_1
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_563_ _563_/A _563_/B _627_/C _563_/D VGND VGND VPWR VPWR _586_/S sky130_fd_sc_hd__or4_1
X_494_ _492_/X _493_/X _492_/X _493_/X VGND VGND VPWR VPWR _494_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_615_ _573_/A _593_/Y _594_/X _595_/X VGND VGND VPWR VPWR _616_/B sky130_fd_sc_hd__o22a_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_546_ _543_/Y _545_/Y _543_/Y _545_/Y VGND VGND VPWR VPWR _546_/X sky130_fd_sc_hd__a2bb2o_1
X_477_ _516_/A _347_/A _544_/A _340_/A VGND VGND VPWR VPWR _479_/A sky130_fd_sc_hd__o22a_1
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_331_ _350_/B VGND VGND VPWR VPWR _436_/A sky130_fd_sc_hd__buf_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_400_ _386_/X _330_/A _392_/Y _391_/B VGND VGND VPWR VPWR _406_/A sky130_fd_sc_hd__a31o_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_529_ _531_/A _531_/C _498_/A VGND VGND VPWR VPWR _529_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_314_ _519_/A _408_/B VGND VGND VPWR VPWR _314_/X sky130_fd_sc_hd__or2_1
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput16 B[7] VGND VGND VPWR VPWR _469_/A sky130_fd_sc_hd__buf_1
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_631_ _631_/A _631_/B VGND VGND VPWR VPWR _631_/Y sky130_fd_sc_hd__nor2_1
X_493_ _457_/X _458_/X _440_/X _459_/X VGND VGND VPWR VPWR _493_/X sky130_fd_sc_hd__o22a_1
X_562_ _563_/A _627_/B _627_/C _584_/A VGND VGND VPWR VPWR _564_/A sky130_fd_sc_hd__o22a_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_476_ _390_/B _469_/X _474_/A _474_/Y _475_/X VGND VGND VPWR VPWR _476_/X sky130_fd_sc_hd__a32o_1
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_614_ _611_/X _613_/X _611_/X _613_/X VGND VGND VPWR VPWR _616_/A sky130_fd_sc_hd__a2bb2o_1
X_545_ _588_/A _584_/A VGND VGND VPWR VPWR _545_/Y sky130_fd_sc_hd__nor2_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _330_/A VGND VGND VPWR VPWR _350_/B sky130_fd_sc_hd__inv_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_459_ _457_/X _458_/X _457_/X _458_/X VGND VGND VPWR VPWR _459_/X sky130_fd_sc_hd__a2bb2o_1
X_528_ _527_/A _527_/B _527_/Y VGND VGND VPWR VPWR _531_/B sky130_fd_sc_hd__a21o_1
XFILLER_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_313_ _313_/A VGND VGND VPWR VPWR _408_/B sky130_fd_sc_hd__buf_1
XFILLER_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_630_ _432_/B _629_/X _432_/B _629_/X VGND VGND VPWR VPWR _630_/X sky130_fd_sc_hd__a2bb2o_1
X_492_ _476_/X _491_/X _476_/X _491_/X VGND VGND VPWR VPWR _492_/X sky130_fd_sc_hd__a2bb2o_1
X_561_ _561_/A VGND VGND VPWR VPWR _627_/C sky130_fd_sc_hd__buf_1
XFILLER_5_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_613_ _588_/A _627_/D _612_/Y _627_/A _586_/S VGND VGND VPWR VPWR _613_/X sky130_fd_sc_hd__o32a_1
X_475_ _475_/A _587_/A VGND VGND VPWR VPWR _475_/X sky130_fd_sc_hd__or2_1
X_544_ _544_/A VGND VGND VPWR VPWR _588_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_458_ _419_/X _420_/X _412_/X _421_/X VGND VGND VPWR VPWR _458_/X sky130_fd_sc_hd__o22a_1
X_527_ _527_/A _527_/B VGND VGND VPWR VPWR _527_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_389_ _442_/D VGND VGND VPWR VPWR _542_/C sky130_fd_sc_hd__buf_1
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_312_ _390_/B VGND VGND VPWR VPWR _313_/A sky130_fd_sc_hd__inv_2
XFILLER_14_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_491_ _489_/X _490_/X _489_/X _490_/X VGND VGND VPWR VPWR _491_/X sky130_fd_sc_hd__a2bb2o_1
X_560_ _563_/B VGND VGND VPWR VPWR _627_/B sky130_fd_sc_hd__buf_1
XFILLER_5_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_474_ _474_/A VGND VGND VPWR VPWR _474_/Y sky130_fd_sc_hd__inv_2
X_612_ _612_/A VGND VGND VPWR VPWR _612_/Y sky130_fd_sc_hd__inv_2
X_543_ _543_/A _543_/B VGND VGND VPWR VPWR _543_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_526_ _504_/X _525_/X _504_/X _525_/X VGND VGND VPWR VPWR _527_/B sky130_fd_sc_hd__a2bb2o_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_457_ _446_/X _456_/X _446_/X _456_/X VGND VGND VPWR VPWR _457_/X sky130_fd_sc_hd__a2bb2o_1
X_388_ _442_/B VGND VGND VPWR VPWR _542_/B sky130_fd_sc_hd__buf_1
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_311_ _447_/B VGND VGND VPWR VPWR _519_/A sky130_fd_sc_hd__buf_1
X_509_ _509_/A VGND VGND VPWR VPWR _509_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_490_ _454_/X _455_/X _446_/X _456_/X VGND VGND VPWR VPWR _490_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_473_ _510_/A _472_/B _471_/Y _471_/A _472_/Y VGND VGND VPWR VPWR _474_/A sky130_fd_sc_hd__o32a_1
X_611_ _591_/A _610_/A _591_/Y _610_/Y VGND VGND VPWR VPWR _611_/X sky130_fd_sc_hd__a22o_1
X_542_ _542_/A _542_/B _542_/C _542_/D VGND VGND VPWR VPWR _543_/B sky130_fd_sc_hd__and4_1
XFILLER_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_387_ _347_/A _313_/A _350_/C _445_/A VGND VGND VPWR VPWR _391_/A sky130_fd_sc_hd__o22a_1
X_525_ _523_/X _524_/X _523_/X _524_/X VGND VGND VPWR VPWR _525_/X sky130_fd_sc_hd__a2bb2o_1
X_456_ _454_/X _455_/X _454_/X _455_/X VGND VGND VPWR VPWR _456_/X sky130_fd_sc_hd__a2bb2o_1
X_310_ _485_/D VGND VGND VPWR VPWR _447_/B sky130_fd_sc_hd__inv_2
X_439_ _437_/X _438_/X _437_/X _438_/X VGND VGND VPWR VPWR _439_/X sky130_fd_sc_hd__a2bb2o_1
X_508_ _539_/A _585_/B _506_/Y _506_/A _507_/Y VGND VGND VPWR VPWR _509_/A sky130_fd_sc_hd__o32a_1
XFILLER_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_472_ _510_/A _472_/B VGND VGND VPWR VPWR _472_/Y sky130_fd_sc_hd__nor2_1
X_610_ _610_/A VGND VGND VPWR VPWR _610_/Y sky130_fd_sc_hd__inv_2
X_541_ _561_/A _347_/A _340_/A _451_/A VGND VGND VPWR VPWR _543_/A sky130_fd_sc_hd__o22a_1
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_524_ _489_/X _490_/X _476_/X _491_/X VGND VGND VPWR VPWR _524_/X sky130_fd_sc_hd__o22a_1
X_455_ _413_/X _418_/X _418_/B VGND VGND VPWR VPWR _455_/X sky130_fd_sc_hd__o21ba_1
X_386_ _386_/A VGND VGND VPWR VPWR _386_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_369_ _342_/X _343_/X _342_/X _343_/X VGND VGND VPWR VPWR _370_/B sky130_fd_sc_hd__a2bb2o_1
X_438_ _475_/A _472_/B VGND VGND VPWR VPWR _438_/X sky130_fd_sc_hd__or2_1
X_507_ _539_/A _585_/B VGND VGND VPWR VPWR _507_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_471_ _471_/A VGND VGND VPWR VPWR _471_/Y sky130_fd_sc_hd__inv_2
X_540_ _410_/C _469_/X _538_/A _538_/Y _539_/X VGND VGND VPWR VPWR _540_/X sky130_fd_sc_hd__a32o_1
XFILLER_20_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_385_ _393_/A VGND VGND VPWR VPWR _386_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_523_ _511_/X _522_/X _511_/X _522_/X VGND VGND VPWR VPWR _523_/X sky130_fd_sc_hd__a2bb2o_1
X_454_ _447_/X _453_/X _447_/X _453_/X VGND VGND VPWR VPWR _454_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_368_ _368_/A _368_/B VGND VGND VPWR VPWR _370_/A sky130_fd_sc_hd__or2_1
X_437_ _408_/X _411_/X _411_/B VGND VGND VPWR VPWR _437_/X sky130_fd_sc_hd__o21ba_1
X_506_ _506_/A VGND VGND VPWR VPWR _506_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_470_ _410_/B _386_/A _444_/Y _443_/B VGND VGND VPWR VPWR _471_/A sky130_fd_sc_hd__a31o_1
X_599_ _599_/A VGND VGND VPWR VPWR _599_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_384_ _375_/X _383_/X _375_/X _383_/X VGND VGND VPWR VPWR _384_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_522_ _520_/X _521_/X _520_/X _521_/X VGND VGND VPWR VPWR _522_/X sky130_fd_sc_hd__a2bb2o_1
X_453_ _381_/C _542_/D _519_/C _449_/A _452_/X VGND VGND VPWR VPWR _453_/X sky130_fd_sc_hd__a32o_1
X_436_ _436_/A _587_/A VGND VGND VPWR VPWR _436_/X sky130_fd_sc_hd__or2_1
X_367_ _631_/A _475_/A _367_/C _631_/B VGND VGND VPWR VPWR _368_/B sky130_fd_sc_hd__or4_1
X_505_ _410_/C _386_/A _480_/Y _479_/B VGND VGND VPWR VPWR _506_/A sky130_fd_sc_hd__a31o_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_419_ _413_/X _418_/X _413_/X _418_/X VGND VGND VPWR VPWR _419_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_598_ _598_/A _598_/B VGND VGND VPWR VPWR _599_/A sky130_fd_sc_hd__or2_1
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_383_ _376_/X _382_/X _376_/X _382_/X VGND VGND VPWR VPWR _383_/X sky130_fd_sc_hd__a2bb2o_1
X_452_ _452_/A _563_/B VGND VGND VPWR VPWR _452_/X sky130_fd_sc_hd__or2_1
X_521_ _486_/X _487_/X _483_/X _488_/X VGND VGND VPWR VPWR _521_/X sky130_fd_sc_hd__o22a_1
XFILLER_16_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_366_ _332_/X _337_/X _332_/X _337_/X VGND VGND VPWR VPWR _368_/A sky130_fd_sc_hd__a2bb2o_1
X_504_ _510_/A _627_/A _471_/Y _474_/Y _475_/X VGND VGND VPWR VPWR _504_/X sky130_fd_sc_hd__o32a_1
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_435_ _570_/B VGND VGND VPWR VPWR _587_/A sky130_fd_sc_hd__buf_1
XFILLER_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_349_ _563_/A _436_/A _350_/C _475_/A VGND VGND VPWR VPWR _351_/A sky130_fd_sc_hd__o22a_1
X_418_ _418_/A _418_/B VGND VGND VPWR VPWR _418_/X sky130_fd_sc_hd__or2_1
XFILLER_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_597_ _574_/X _575_/X _559_/X _576_/X VGND VGND VPWR VPWR _598_/B sky130_fd_sc_hd__o22a_1
XFILLER_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_520_ _518_/X _519_/X _518_/X _519_/X VGND VGND VPWR VPWR _520_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_382_ _382_/A _382_/B VGND VGND VPWR VPWR _382_/X sky130_fd_sc_hd__or2_1
X_451_ _451_/A VGND VGND VPWR VPWR _563_/B sky130_fd_sc_hd__buf_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_365_ _363_/A _363_/B _629_/A VGND VGND VPWR VPWR _371_/A sky130_fd_sc_hd__a21o_1
X_503_ _503_/A VGND VGND VPWR VPWR _627_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_434_ _469_/A VGND VGND VPWR VPWR _570_/B sky130_fd_sc_hd__inv_2
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_348_ _408_/B VGND VGND VPWR VPWR _475_/A sky130_fd_sc_hd__buf_1
X_417_ _417_/A _513_/A _542_/A _417_/D VGND VGND VPWR VPWR _418_/B sky130_fd_sc_hd__and4_1
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_596_ _594_/X _595_/X _594_/X _595_/X VGND VGND VPWR VPWR _598_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_381_ _485_/A _381_/B _381_/C _513_/A VGND VGND VPWR VPWR _382_/B sky130_fd_sc_hd__and4_1
X_450_ _542_/D VGND VGND VPWR VPWR _451_/A sky130_fd_sc_hd__inv_2
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_579_ _580_/A _580_/B VGND VGND VPWR VPWR _579_/X sky130_fd_sc_hd__and2_1
X_433_ _431_/X _432_/X _431_/X _432_/X VGND VGND VPWR VPWR _433_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_502_ _492_/X _493_/X _468_/X _494_/X VGND VGND VPWR VPWR _527_/A sky130_fd_sc_hd__o22a_1
X_364_ _430_/A VGND VGND VPWR VPWR _629_/A sky130_fd_sc_hd__inv_2
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_347_ _347_/A VGND VGND VPWR VPWR _563_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_416_ _448_/B _378_/A _561_/A _452_/A VGND VGND VPWR VPWR _418_/A sky130_fd_sc_hd__o22a_1
XFILLER_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_595_ _588_/A _627_/A _566_/Y _569_/Y _570_/X VGND VGND VPWR VPWR _595_/X sky130_fd_sc_hd__o32a_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput30 _467_/Y VGND VGND VPWR VPWR M[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_380_ _380_/A VGND VGND VPWR VPWR _513_/A sky130_fd_sc_hd__buf_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_578_ _549_/X _550_/X _533_/X _551_/X VGND VGND VPWR VPWR _580_/B sky130_fd_sc_hd__o22a_1
.ends


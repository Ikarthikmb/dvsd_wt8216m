magic
tech sky130A
magscale 1 2
timestamp 1629484573
<< checkpaint >>
rect -3932 -3932 21516 23660
<< locali >>
rect 16589 10251 16623 12733
rect 16681 10659 16715 11645
rect 4813 6103 4847 6273
rect 12817 5151 12851 5253
rect 16681 5151 16715 10625
rect 13921 2431 13955 2601
<< viali >>
rect 2605 17289 2639 17323
rect 12633 17289 12667 17323
rect 1869 17221 1903 17255
rect 4169 17221 4203 17255
rect 8033 17221 8067 17255
rect 9965 17221 9999 17255
rect 10885 17221 10919 17255
rect 2697 17153 2731 17187
rect 4353 17153 4387 17187
rect 5089 17153 5123 17187
rect 5641 17153 5675 17187
rect 6377 17153 6411 17187
rect 8217 17153 8251 17187
rect 9229 17153 9263 17187
rect 9413 17153 9447 17187
rect 10149 17153 10183 17187
rect 10793 17153 10827 17187
rect 11713 17153 11747 17187
rect 11805 17153 11839 17187
rect 12081 17153 12115 17187
rect 12725 17153 12759 17187
rect 13461 17153 13495 17187
rect 14289 17153 14323 17187
rect 15025 17153 15059 17187
rect 15577 17153 15611 17187
rect 2053 17085 2087 17119
rect 6653 17085 6687 17119
rect 4905 17017 4939 17051
rect 14841 17017 14875 17051
rect 15761 17017 15795 17051
rect 5733 16949 5767 16983
rect 9045 16949 9079 16983
rect 10333 16949 10367 16983
rect 11529 16949 11563 16983
rect 11989 16949 12023 16983
rect 13277 16949 13311 16983
rect 14105 16949 14139 16983
rect 2329 16745 2363 16779
rect 8125 16745 8159 16779
rect 12173 16745 12207 16779
rect 14657 16745 14691 16779
rect 4077 16677 4111 16711
rect 4813 16677 4847 16711
rect 14197 16677 14231 16711
rect 2053 16609 2087 16643
rect 3801 16609 3835 16643
rect 4353 16609 4387 16643
rect 6285 16609 6319 16643
rect 6929 16609 6963 16643
rect 7389 16609 7423 16643
rect 9045 16609 9079 16643
rect 9873 16609 9907 16643
rect 10333 16609 10367 16643
rect 11529 16609 11563 16643
rect 11989 16609 12023 16643
rect 13093 16609 13127 16643
rect 13553 16609 13587 16643
rect 2237 16541 2271 16575
rect 2605 16541 2639 16575
rect 3939 16541 3973 16575
rect 4169 16541 4203 16575
rect 4997 16541 5031 16575
rect 5365 16541 5399 16575
rect 5825 16541 5859 16575
rect 6101 16541 6135 16575
rect 7021 16541 7055 16575
rect 7297 16541 7331 16575
rect 8125 16541 8159 16575
rect 8401 16541 8435 16575
rect 9413 16541 9447 16575
rect 9965 16541 9999 16575
rect 10241 16541 10275 16575
rect 11621 16541 11655 16575
rect 11897 16541 11931 16575
rect 13185 16541 13219 16575
rect 14105 16541 14139 16575
rect 14381 16541 14415 16575
rect 14473 16541 14507 16575
rect 5089 16473 5123 16507
rect 5181 16473 5215 16507
rect 9229 16473 9263 16507
rect 13461 16473 13495 16507
rect 15209 16473 15243 16507
rect 15393 16473 15427 16507
rect 2513 16405 2547 16439
rect 5917 16405 5951 16439
rect 7573 16405 7607 16439
rect 8309 16405 8343 16439
rect 10517 16405 10551 16439
rect 12909 16405 12943 16439
rect 15577 16405 15611 16439
rect 4905 16201 4939 16235
rect 5457 16201 5491 16235
rect 8217 16201 8251 16235
rect 9229 16201 9263 16235
rect 11529 16201 11563 16235
rect 15393 16201 15427 16235
rect 5641 16133 5675 16167
rect 9413 16133 9447 16167
rect 10149 16133 10183 16167
rect 10517 16133 10551 16167
rect 13553 16133 13587 16167
rect 15301 16133 15335 16167
rect 3709 16065 3743 16099
rect 3801 16065 3835 16099
rect 4077 16065 4111 16099
rect 4813 16065 4847 16099
rect 5825 16065 5859 16099
rect 6745 16065 6779 16099
rect 6837 16065 6871 16099
rect 7113 16065 7147 16099
rect 7941 16065 7975 16099
rect 9597 16065 9631 16099
rect 10333 16065 10367 16099
rect 10609 16065 10643 16099
rect 11805 16065 11839 16099
rect 12081 16065 12115 16099
rect 13277 16065 13311 16099
rect 13645 16065 13679 16099
rect 14565 16065 14599 16099
rect 15209 16065 15243 16099
rect 7757 15997 7791 16031
rect 8309 15997 8343 16031
rect 11713 15997 11747 16031
rect 12173 15997 12207 16031
rect 13185 15997 13219 16031
rect 15669 15997 15703 16031
rect 6561 15929 6595 15963
rect 7021 15929 7055 15963
rect 13001 15929 13035 15963
rect 14749 15929 14783 15963
rect 3525 15861 3559 15895
rect 3985 15861 4019 15895
rect 8033 15861 8067 15895
rect 1593 15657 1627 15691
rect 2513 15657 2547 15691
rect 9965 15657 9999 15691
rect 13001 15657 13035 15691
rect 13185 15657 13219 15691
rect 15209 15657 15243 15691
rect 1685 15589 1719 15623
rect 2697 15521 2731 15555
rect 3801 15521 3835 15555
rect 1777 15453 1811 15487
rect 2421 15453 2455 15487
rect 9873 15453 9907 15487
rect 10517 15453 10551 15487
rect 10885 15453 10919 15487
rect 11621 15453 11655 15487
rect 12081 15453 12115 15487
rect 12725 15453 12759 15487
rect 14657 15453 14691 15487
rect 14933 15453 14967 15487
rect 15025 15453 15059 15487
rect 1501 15385 1535 15419
rect 3985 15385 4019 15419
rect 4169 15385 4203 15419
rect 10701 15385 10735 15419
rect 14565 15385 14599 15419
rect 2697 15317 2731 15351
rect 11437 15317 11471 15351
rect 12265 15317 12299 15351
rect 3801 15113 3835 15147
rect 6469 15113 6503 15147
rect 7849 15113 7883 15147
rect 12173 15113 12207 15147
rect 13645 15113 13679 15147
rect 15301 15113 15335 15147
rect 5549 15045 5583 15079
rect 7021 15045 7055 15079
rect 2145 14977 2179 15011
rect 2421 14977 2455 15011
rect 3341 14977 3375 15011
rect 3985 14977 4019 15011
rect 4077 14977 4111 15011
rect 5181 14977 5215 15011
rect 6745 14977 6779 15011
rect 8125 14977 8159 15011
rect 8401 14977 8435 15011
rect 11529 14977 11563 15011
rect 11897 14977 11931 15011
rect 12633 14977 12667 15011
rect 13829 14977 13863 15011
rect 13921 14977 13955 15011
rect 14197 14977 14231 15011
rect 14657 14977 14691 15011
rect 15025 14977 15059 15011
rect 2053 14909 2087 14943
rect 2513 14909 2547 14943
rect 4353 14909 4387 14943
rect 4445 14909 4479 14943
rect 5089 14909 5123 14943
rect 5457 14909 5491 14943
rect 6653 14909 6687 14943
rect 7113 14909 7147 14943
rect 8033 14909 8067 14943
rect 8493 14909 8527 14943
rect 11621 14909 11655 14943
rect 11989 14909 12023 14943
rect 14749 14909 14783 14943
rect 15117 14909 15151 14943
rect 4905 14841 4939 14875
rect 14105 14841 14139 14875
rect 2697 14773 2731 14807
rect 3249 14773 3283 14807
rect 12817 14773 12851 14807
rect 2789 14569 2823 14603
rect 4261 14569 4295 14603
rect 4721 14569 4755 14603
rect 7113 14569 7147 14603
rect 7573 14569 7607 14603
rect 8953 14569 8987 14603
rect 11345 14569 11379 14603
rect 12357 14569 12391 14603
rect 14841 14569 14875 14603
rect 15393 14569 15427 14603
rect 11805 14433 11839 14467
rect 14289 14433 14323 14467
rect 1961 14365 1995 14399
rect 2973 14365 3007 14399
rect 3157 14365 3191 14399
rect 3249 14365 3283 14399
rect 4445 14365 4479 14399
rect 4537 14365 4571 14399
rect 4813 14365 4847 14399
rect 7297 14365 7331 14399
rect 7389 14365 7423 14399
rect 7665 14365 7699 14399
rect 8125 14365 8159 14399
rect 8309 14365 8343 14399
rect 9137 14365 9171 14399
rect 9229 14365 9263 14399
rect 9505 14365 9539 14399
rect 10701 14365 10735 14399
rect 10885 14365 10919 14399
rect 11529 14365 11563 14399
rect 11621 14365 11655 14399
rect 11897 14365 11931 14399
rect 12541 14365 12575 14399
rect 12633 14365 12667 14399
rect 12909 14365 12943 14399
rect 14565 14365 14599 14399
rect 14657 14365 14691 14399
rect 15577 14365 15611 14399
rect 9597 14297 9631 14331
rect 13001 14297 13035 14331
rect 14197 14297 14231 14331
rect 15761 14297 15795 14331
rect 1777 14229 1811 14263
rect 8217 14229 8251 14263
rect 10793 14229 10827 14263
rect 2237 14025 2271 14059
rect 7205 14025 7239 14059
rect 8033 14025 8067 14059
rect 11529 14025 11563 14059
rect 13737 14025 13771 14059
rect 15577 14025 15611 14059
rect 1501 13957 1535 13991
rect 9965 13957 9999 13991
rect 11897 13957 11931 13991
rect 1593 13889 1627 13923
rect 2234 13889 2268 13923
rect 2697 13889 2731 13923
rect 3525 13889 3559 13923
rect 3617 13889 3651 13923
rect 3893 13889 3927 13923
rect 5089 13889 5123 13923
rect 5181 13889 5215 13923
rect 5457 13889 5491 13923
rect 7389 13889 7423 13923
rect 7481 13889 7515 13923
rect 7941 13889 7975 13923
rect 8125 13889 8159 13923
rect 9597 13889 9631 13923
rect 9873 13889 9907 13923
rect 10977 13889 11011 13923
rect 11713 13889 11747 13923
rect 11805 13889 11839 13923
rect 12015 13889 12049 13923
rect 12817 13889 12851 13923
rect 13921 13889 13955 13923
rect 14197 13889 14231 13923
rect 14381 13889 14415 13923
rect 15301 13889 15335 13923
rect 15669 13889 15703 13923
rect 15761 13889 15795 13923
rect 3341 13821 3375 13855
rect 7205 13821 7239 13855
rect 9505 13821 9539 13855
rect 10885 13821 10919 13855
rect 12173 13821 12207 13855
rect 2053 13685 2087 13719
rect 2605 13685 2639 13719
rect 3801 13685 3835 13719
rect 4905 13685 4939 13719
rect 5365 13685 5399 13719
rect 9321 13685 9355 13719
rect 12725 13685 12759 13719
rect 2145 13481 2179 13515
rect 3065 13481 3099 13515
rect 3801 13481 3835 13515
rect 4997 13481 5031 13515
rect 10977 13481 11011 13515
rect 12357 13481 12391 13515
rect 13553 13481 13587 13515
rect 14473 13481 14507 13515
rect 9413 13413 9447 13447
rect 11161 13345 11195 13379
rect 11253 13345 11287 13379
rect 2329 13277 2363 13311
rect 2605 13277 2639 13311
rect 3065 13277 3099 13311
rect 3249 13277 3283 13311
rect 3985 13277 4019 13311
rect 4077 13277 4111 13311
rect 4353 13277 4387 13311
rect 5181 13277 5215 13311
rect 5273 13277 5307 13311
rect 5549 13277 5583 13311
rect 7665 13277 7699 13311
rect 9137 13277 9171 13311
rect 9229 13277 9263 13311
rect 9505 13277 9539 13311
rect 10333 13277 10367 13311
rect 11345 13277 11379 13311
rect 11437 13277 11471 13311
rect 2513 13209 2547 13243
rect 4445 13209 4479 13243
rect 5641 13209 5675 13243
rect 7849 13209 7883 13243
rect 11989 13209 12023 13243
rect 12173 13209 12207 13243
rect 13185 13209 13219 13243
rect 13369 13209 13403 13243
rect 14105 13209 14139 13243
rect 14289 13209 14323 13243
rect 14933 13209 14967 13243
rect 15117 13209 15151 13243
rect 7481 13141 7515 13175
rect 8953 13141 8987 13175
rect 10425 13141 10459 13175
rect 15301 13141 15335 13175
rect 3433 12937 3467 12971
rect 5181 12937 5215 12971
rect 6561 12937 6595 12971
rect 9413 12937 9447 12971
rect 11897 12937 11931 12971
rect 13185 12937 13219 12971
rect 14381 12937 14415 12971
rect 15025 12937 15059 12971
rect 1961 12869 1995 12903
rect 4077 12869 4111 12903
rect 5733 12869 5767 12903
rect 7205 12869 7239 12903
rect 10701 12869 10735 12903
rect 14013 12869 14047 12903
rect 2513 12801 2547 12835
rect 2697 12801 2731 12835
rect 3617 12801 3651 12835
rect 3709 12801 3743 12835
rect 3985 12801 4019 12835
rect 5457 12801 5491 12835
rect 5825 12801 5859 12835
rect 6745 12801 6779 12835
rect 6837 12801 6871 12835
rect 7941 12801 7975 12835
rect 8217 12801 8251 12835
rect 8769 12801 8803 12835
rect 9689 12801 9723 12835
rect 9965 12801 9999 12835
rect 10885 12801 10919 12835
rect 11529 12801 11563 12835
rect 11713 12801 11747 12835
rect 12633 12801 12667 12835
rect 12909 12801 12943 12835
rect 13001 12801 13035 12835
rect 14197 12801 14231 12835
rect 15209 12801 15243 12835
rect 15485 12801 15519 12835
rect 15669 12801 15703 12835
rect 5365 12733 5399 12767
rect 7113 12733 7147 12767
rect 7849 12733 7883 12767
rect 8309 12733 8343 12767
rect 9597 12733 9631 12767
rect 10057 12733 10091 12767
rect 10517 12733 10551 12767
rect 16589 12733 16623 12767
rect 12725 12665 12759 12699
rect 1869 12597 1903 12631
rect 2513 12597 2547 12631
rect 7665 12597 7699 12631
rect 8953 12597 8987 12631
rect 1593 12393 1627 12427
rect 7205 12393 7239 12427
rect 11621 12393 11655 12427
rect 12265 12393 12299 12427
rect 12725 12393 12759 12427
rect 14657 12393 14691 12427
rect 15761 12393 15795 12427
rect 1869 12325 1903 12359
rect 1961 12257 1995 12291
rect 2789 12257 2823 12291
rect 7665 12257 7699 12291
rect 9229 12257 9263 12291
rect 10885 12257 10919 12291
rect 12633 12257 12667 12291
rect 14197 12257 14231 12291
rect 1777 12189 1811 12223
rect 2053 12189 2087 12223
rect 2237 12189 2271 12223
rect 2881 12189 2915 12223
rect 7389 12189 7423 12223
rect 7481 12189 7515 12223
rect 7757 12189 7791 12223
rect 8217 12189 8251 12223
rect 9413 12189 9447 12223
rect 9689 12189 9723 12223
rect 9873 12189 9907 12223
rect 11161 12189 11195 12223
rect 11805 12189 11839 12223
rect 12449 12189 12483 12223
rect 13185 12189 13219 12223
rect 14105 12189 14139 12223
rect 14381 12189 14415 12223
rect 14473 12189 14507 12223
rect 15209 12189 15243 12223
rect 15485 12189 15519 12223
rect 15577 12189 15611 12223
rect 12725 12121 12759 12155
rect 13369 12121 13403 12155
rect 13553 12121 13587 12155
rect 15117 12121 15151 12155
rect 8401 12053 8435 12087
rect 2881 11849 2915 11883
rect 3985 11849 4019 11883
rect 5181 11849 5215 11883
rect 8033 11849 8067 11883
rect 9689 11849 9723 11883
rect 12173 11849 12207 11883
rect 14289 11849 14323 11883
rect 15669 11849 15703 11883
rect 5825 11781 5859 11815
rect 8401 11781 8435 11815
rect 9321 11781 9355 11815
rect 15209 11781 15243 11815
rect 2053 11713 2087 11747
rect 2237 11713 2271 11747
rect 3157 11713 3191 11747
rect 4169 11713 4203 11747
rect 4261 11713 4295 11747
rect 5365 11713 5399 11747
rect 5457 11713 5491 11747
rect 7113 11713 7147 11747
rect 7297 11713 7331 11747
rect 7573 11713 7607 11747
rect 8217 11713 8251 11747
rect 9505 11713 9539 11747
rect 10977 11713 11011 11747
rect 11621 11713 11655 11747
rect 11897 11713 11931 11747
rect 11989 11713 12023 11747
rect 12817 11713 12851 11747
rect 13737 11713 13771 11747
rect 14013 11713 14047 11747
rect 14105 11713 14139 11747
rect 15485 11713 15519 11747
rect 2145 11645 2179 11679
rect 2329 11645 2363 11679
rect 3065 11645 3099 11679
rect 3433 11645 3467 11679
rect 3525 11645 3559 11679
rect 4537 11645 4571 11679
rect 4629 11645 4663 11679
rect 5733 11645 5767 11679
rect 7389 11645 7423 11679
rect 10701 11645 10735 11679
rect 11713 11645 11747 11679
rect 12725 11645 12759 11679
rect 15393 11645 15427 11679
rect 6929 11577 6963 11611
rect 7205 11577 7239 11611
rect 13829 11577 13863 11611
rect 1869 11509 1903 11543
rect 15209 11509 15243 11543
rect 3893 11305 3927 11339
rect 11529 11305 11563 11339
rect 15393 11305 15427 11339
rect 13369 11237 13403 11271
rect 1685 11169 1719 11203
rect 2145 11169 2179 11203
rect 3157 11169 3191 11203
rect 7573 11169 7607 11203
rect 8401 11169 8435 11203
rect 9689 11169 9723 11203
rect 11989 11169 12023 11203
rect 12633 11169 12667 11203
rect 14381 11169 14415 11203
rect 1869 11101 1903 11135
rect 1961 11101 1995 11135
rect 2053 11101 2087 11135
rect 2881 11101 2915 11135
rect 2973 11101 3007 11135
rect 3249 11101 3283 11135
rect 4077 11101 4111 11135
rect 4169 11101 4203 11135
rect 4445 11101 4479 11135
rect 6285 11101 6319 11135
rect 6469 11101 6503 11135
rect 7114 11079 7148 11113
rect 7297 11101 7331 11135
rect 8225 11101 8259 11135
rect 9597 11101 9631 11135
rect 9781 11101 9815 11135
rect 9873 11101 9907 11135
rect 10609 11101 10643 11135
rect 11713 11101 11747 11135
rect 11805 11101 11839 11135
rect 12081 11101 12115 11135
rect 12725 11101 12759 11135
rect 13185 11101 13219 11135
rect 14105 11101 14139 11135
rect 15577 11101 15611 11135
rect 15761 11101 15795 11135
rect 2697 11033 2731 11067
rect 4537 11033 4571 11067
rect 6377 11033 6411 11067
rect 7205 11033 7239 11067
rect 7415 11033 7449 11067
rect 8033 11033 8067 11067
rect 6929 10965 6963 10999
rect 9413 10965 9447 10999
rect 10425 10965 10459 10999
rect 2789 10761 2823 10795
rect 3893 10761 3927 10795
rect 4905 10761 4939 10795
rect 6561 10761 6595 10795
rect 10701 10761 10735 10795
rect 10977 10761 11011 10795
rect 13277 10761 13311 10795
rect 15485 10761 15519 10795
rect 9597 10693 9631 10727
rect 9827 10693 9861 10727
rect 11529 10693 11563 10727
rect 11713 10693 11747 10727
rect 12909 10693 12943 10727
rect 2145 10625 2179 10659
rect 2237 10625 2271 10659
rect 2697 10625 2731 10659
rect 4077 10625 4111 10659
rect 4169 10625 4203 10659
rect 4445 10625 4479 10659
rect 5181 10625 5215 10659
rect 5457 10625 5491 10659
rect 6653 10625 6687 10659
rect 7297 10625 7331 10659
rect 9505 10625 9539 10659
rect 9689 10625 9723 10659
rect 10609 10625 10643 10659
rect 10793 10625 10827 10659
rect 11897 10625 11931 10659
rect 12725 10625 12759 10659
rect 13001 10625 13035 10659
rect 13093 10625 13127 10659
rect 13921 10625 13955 10659
rect 14933 10625 14967 10659
rect 15209 10625 15243 10659
rect 15301 10625 15335 10659
rect 1961 10557 1995 10591
rect 4353 10557 4387 10591
rect 5089 10557 5123 10591
rect 5549 10557 5583 10591
rect 7757 10557 7791 10591
rect 8033 10557 8067 10591
rect 9965 10557 9999 10591
rect 9321 10489 9355 10523
rect 10425 10489 10459 10523
rect 13737 10489 13771 10523
rect 15025 10489 15059 10523
rect 2053 10421 2087 10455
rect 7205 10421 7239 10455
rect 2605 10217 2639 10251
rect 5457 10217 5491 10251
rect 7757 10217 7791 10251
rect 9781 10217 9815 10251
rect 12081 10217 12115 10251
rect 13277 10217 13311 10251
rect 16589 10217 16623 10251
rect 16681 11645 16715 11679
rect 16681 10625 16715 10659
rect 1501 10081 1535 10115
rect 1961 10081 1995 10115
rect 2789 10081 2823 10115
rect 5917 10081 5951 10115
rect 8033 10081 8067 10115
rect 8217 10081 8251 10115
rect 10333 10081 10367 10115
rect 11161 10081 11195 10115
rect 15393 10081 15427 10115
rect 1593 10013 1627 10047
rect 1869 10013 1903 10047
rect 2881 10013 2915 10047
rect 3249 10013 3283 10047
rect 3801 10013 3835 10047
rect 5641 10013 5675 10047
rect 5733 10013 5767 10047
rect 6009 10013 6043 10047
rect 7113 10013 7147 10047
rect 7941 10013 7975 10047
rect 8134 10013 8168 10047
rect 8401 10013 8435 10047
rect 8953 10013 8987 10047
rect 10149 10013 10183 10047
rect 13093 10013 13127 10047
rect 14105 10013 14139 10047
rect 15117 10013 15151 10047
rect 3985 9945 4019 9979
rect 6929 9945 6963 9979
rect 10793 9945 10827 9979
rect 10977 9945 11011 9979
rect 11989 9945 12023 9979
rect 12725 9945 12759 9979
rect 14289 9945 14323 9979
rect 2145 9877 2179 9911
rect 4169 9877 4203 9911
rect 7297 9877 7331 9911
rect 9137 9877 9171 9911
rect 9965 9877 9999 9911
rect 10057 9877 10091 9911
rect 12909 9877 12943 9911
rect 13001 9877 13035 9911
rect 14473 9877 14507 9911
rect 1869 9673 1903 9707
rect 8493 9673 8527 9707
rect 9689 9673 9723 9707
rect 5733 9605 5767 9639
rect 12173 9605 12207 9639
rect 14657 9605 14691 9639
rect 2144 9537 2178 9571
rect 2237 9537 2271 9571
rect 2881 9537 2915 9571
rect 2973 9537 3007 9571
rect 5457 9537 5491 9571
rect 7297 9537 7331 9571
rect 7573 9537 7607 9571
rect 7757 9537 7791 9571
rect 8585 9537 8619 9571
rect 9045 9537 9079 9571
rect 9873 9537 9907 9571
rect 9965 9537 9999 9571
rect 10057 9537 10091 9571
rect 10793 9537 10827 9571
rect 10885 9537 10919 9571
rect 11805 9537 11839 9571
rect 13093 9537 13127 9571
rect 13829 9537 13863 9571
rect 14105 9537 14139 9571
rect 14841 9537 14875 9571
rect 15117 9537 15151 9571
rect 15301 9537 15335 9571
rect 2697 9469 2731 9503
rect 5365 9469 5399 9503
rect 5825 9469 5859 9503
rect 7481 9469 7515 9503
rect 13737 9469 13771 9503
rect 14197 9469 14231 9503
rect 2789 9401 2823 9435
rect 7389 9401 7423 9435
rect 10241 9401 10275 9435
rect 13553 9401 13587 9435
rect 5181 9333 5215 9367
rect 7113 9333 7147 9367
rect 9229 9333 9263 9367
rect 12909 9333 12943 9367
rect 2145 9129 2179 9163
rect 3893 9129 3927 9163
rect 11161 9129 11195 9163
rect 11621 9129 11655 9163
rect 13553 9129 13587 9163
rect 14105 9129 14139 9163
rect 4077 8993 4111 9027
rect 4537 8993 4571 9027
rect 7297 8993 7331 9027
rect 7941 8993 7975 9027
rect 9229 8993 9263 9027
rect 10609 8993 10643 9027
rect 12449 8993 12483 9027
rect 2789 8925 2823 8959
rect 4169 8925 4203 8959
rect 6837 8925 6871 8959
rect 7481 8925 7515 8959
rect 7665 8925 7699 8959
rect 8953 8925 8987 8959
rect 10517 8925 10551 8959
rect 11345 8925 11379 8959
rect 11437 8925 11471 8959
rect 11713 8925 11747 8959
rect 13369 8925 13403 8959
rect 14289 8925 14323 8959
rect 14565 8925 14599 8959
rect 14749 8925 14783 8959
rect 1777 8857 1811 8891
rect 1961 8857 1995 8891
rect 4445 8857 4479 8891
rect 6745 8857 6779 8891
rect 7573 8857 7607 8891
rect 7783 8857 7817 8891
rect 12265 8857 12299 8891
rect 13185 8857 13219 8891
rect 15485 8857 15519 8891
rect 15669 8857 15703 8891
rect 2697 8789 2731 8823
rect 1685 8585 1719 8619
rect 3157 8585 3191 8619
rect 5181 8585 5215 8619
rect 8033 8585 8067 8619
rect 10149 8585 10183 8619
rect 13093 8585 13127 8619
rect 13277 8585 13311 8619
rect 13461 8585 13495 8619
rect 6929 8517 6963 8551
rect 9413 8517 9447 8551
rect 14105 8517 14139 8551
rect 1869 8449 1903 8483
rect 2605 8449 2639 8483
rect 2881 8449 2915 8483
rect 2973 8449 3007 8483
rect 4353 8449 4387 8483
rect 4629 8449 4663 8483
rect 5457 8449 5491 8483
rect 8217 8449 8251 8483
rect 8493 8449 8527 8483
rect 8677 8449 8711 8483
rect 9321 8449 9355 8483
rect 9965 8449 9999 8483
rect 10241 8449 10275 8483
rect 10333 8449 10367 8483
rect 11805 8449 11839 8483
rect 13185 8449 13219 8483
rect 14289 8449 14323 8483
rect 15209 8449 15243 8483
rect 15485 8449 15519 8483
rect 2053 8381 2087 8415
rect 2513 8381 2547 8415
rect 4261 8381 4295 8415
rect 4721 8381 4755 8415
rect 5365 8381 5399 8415
rect 5733 8381 5767 8415
rect 5825 8381 5859 8415
rect 8401 8381 8435 8415
rect 12081 8381 12115 8415
rect 14473 8381 14507 8415
rect 15117 8381 15151 8415
rect 15577 8381 15611 8415
rect 4077 8313 4111 8347
rect 8309 8313 8343 8347
rect 12909 8313 12943 8347
rect 14933 8313 14967 8347
rect 7021 8245 7055 8279
rect 10517 8245 10551 8279
rect 2513 8041 2547 8075
rect 5549 8041 5583 8075
rect 6653 8041 6687 8075
rect 8309 8041 8343 8075
rect 12357 8041 12391 8075
rect 14105 8041 14139 8075
rect 14565 8041 14599 8075
rect 15485 8041 15519 8075
rect 6193 7973 6227 8007
rect 10425 7973 10459 8007
rect 4629 7905 4663 7939
rect 10701 7905 10735 7939
rect 10793 7905 10827 7939
rect 13001 7905 13035 7939
rect 2697 7837 2731 7871
rect 2789 7837 2823 7871
rect 3065 7837 3099 7871
rect 4169 7837 4203 7871
rect 4353 7837 4387 7871
rect 4445 7837 4479 7871
rect 4721 7837 4755 7871
rect 5365 7837 5399 7871
rect 6009 7837 6043 7871
rect 6653 7837 6687 7871
rect 6837 7837 6871 7871
rect 7481 7837 7515 7871
rect 8401 7837 8435 7871
rect 9505 7837 9539 7871
rect 9689 7837 9723 7871
rect 9965 7837 9999 7871
rect 10609 7837 10643 7871
rect 10885 7837 10919 7871
rect 12449 7837 12483 7871
rect 13277 7837 13311 7871
rect 14289 7837 14323 7871
rect 14381 7837 14415 7871
rect 14657 7837 14691 7871
rect 3157 7769 3191 7803
rect 7665 7769 7699 7803
rect 9597 7769 9631 7803
rect 9827 7769 9861 7803
rect 11437 7769 11471 7803
rect 11621 7769 11655 7803
rect 11805 7769 11839 7803
rect 13553 7769 13587 7803
rect 15117 7769 15151 7803
rect 15301 7769 15335 7803
rect 7297 7701 7331 7735
rect 9321 7701 9355 7735
rect 13185 7701 13219 7735
rect 13369 7701 13403 7735
rect 2237 7497 2271 7531
rect 4169 7497 4203 7531
rect 5273 7497 5307 7531
rect 8769 7497 8803 7531
rect 9965 7497 9999 7531
rect 15117 7497 15151 7531
rect 7021 7429 7055 7463
rect 7757 7429 7791 7463
rect 7849 7429 7883 7463
rect 10701 7429 10735 7463
rect 11529 7429 11563 7463
rect 2421 7361 2455 7395
rect 2513 7361 2547 7395
rect 2789 7361 2823 7395
rect 3985 7361 4019 7395
rect 4629 7361 4663 7395
rect 5457 7361 5491 7395
rect 5549 7361 5583 7395
rect 5825 7361 5859 7395
rect 6561 7361 6595 7395
rect 6653 7361 6687 7395
rect 7665 7361 7699 7395
rect 7987 7361 8021 7395
rect 8585 7361 8619 7395
rect 9413 7361 9447 7395
rect 10057 7361 10091 7395
rect 10517 7361 10551 7395
rect 10885 7361 10919 7395
rect 11713 7361 11747 7395
rect 11805 7361 11839 7395
rect 12081 7361 12115 7395
rect 12541 7361 12575 7395
rect 12725 7361 12759 7395
rect 13829 7361 13863 7395
rect 14565 7361 14599 7395
rect 14841 7361 14875 7395
rect 14933 7361 14967 7395
rect 15577 7361 15611 7395
rect 2697 7293 2731 7327
rect 6929 7293 6963 7327
rect 8125 7293 8159 7327
rect 14657 7293 14691 7327
rect 4813 7225 4847 7259
rect 6377 7225 6411 7259
rect 5733 7157 5767 7191
rect 7481 7157 7515 7191
rect 9229 7157 9263 7191
rect 11989 7157 12023 7191
rect 12909 7157 12943 7191
rect 13645 7157 13679 7191
rect 15669 7157 15703 7191
rect 2421 6953 2455 6987
rect 3801 6953 3835 6987
rect 12817 6953 12851 6987
rect 8033 6885 8067 6919
rect 2605 6817 2639 6851
rect 3985 6817 4019 6851
rect 4445 6817 4479 6851
rect 6101 6817 6135 6851
rect 7113 6817 7147 6851
rect 8125 6817 8159 6851
rect 10011 6817 10045 6851
rect 11345 6817 11379 6851
rect 13461 6817 13495 6851
rect 15669 6817 15703 6851
rect 1409 6749 1443 6783
rect 2697 6749 2731 6783
rect 2973 6749 3007 6783
rect 4077 6749 4111 6783
rect 4353 6749 4387 6783
rect 5365 6749 5399 6783
rect 5549 6749 5583 6783
rect 6193 6749 6227 6783
rect 6837 6749 6871 6783
rect 6929 6749 6963 6783
rect 7021 6749 7055 6783
rect 7297 6749 7331 6783
rect 7941 6749 7975 6783
rect 8217 6749 8251 6783
rect 8401 6749 8435 6783
rect 9505 6749 9539 6783
rect 10241 6749 10275 6783
rect 11713 6749 11747 6783
rect 11805 6749 11839 6783
rect 11989 6749 12023 6783
rect 13001 6749 13035 6783
rect 13093 6749 13127 6783
rect 14197 6749 14231 6783
rect 14565 6749 14599 6783
rect 15209 6749 15243 6783
rect 15301 6749 15335 6783
rect 15577 6749 15611 6783
rect 3065 6681 3099 6715
rect 11483 6681 11517 6715
rect 11608 6681 11642 6715
rect 13369 6681 13403 6715
rect 14381 6681 14415 6715
rect 1593 6613 1627 6647
rect 5457 6613 5491 6647
rect 6653 6613 6687 6647
rect 7757 6613 7791 6647
rect 9321 6613 9355 6647
rect 15025 6613 15059 6647
rect 3249 6409 3283 6443
rect 4905 6409 4939 6443
rect 8125 6409 8159 6443
rect 8769 6409 8803 6443
rect 12081 6409 12115 6443
rect 9413 6341 9447 6375
rect 12265 6341 12299 6375
rect 14749 6341 14783 6375
rect 1685 6273 1719 6307
rect 3433 6273 3467 6307
rect 3525 6273 3559 6307
rect 4813 6273 4847 6307
rect 5181 6273 5215 6307
rect 6561 6273 6595 6307
rect 7205 6273 7239 6307
rect 7389 6273 7423 6307
rect 8033 6273 8067 6307
rect 8217 6273 8251 6307
rect 8861 6273 8895 6307
rect 9505 6273 9539 6307
rect 10241 6273 10275 6307
rect 10425 6273 10459 6307
rect 12449 6273 12483 6307
rect 13093 6273 13127 6307
rect 13369 6273 13403 6307
rect 13553 6273 13587 6307
rect 14105 6273 14139 6307
rect 14933 6273 14967 6307
rect 15209 6273 15243 6307
rect 15393 6273 15427 6307
rect 1409 6205 1443 6239
rect 3801 6205 3835 6239
rect 3893 6205 3927 6239
rect 5089 6205 5123 6239
rect 5457 6205 5491 6239
rect 5549 6205 5583 6239
rect 6469 6205 6503 6239
rect 7021 6205 7055 6239
rect 9965 6205 9999 6239
rect 10149 6205 10183 6239
rect 10333 6205 10367 6239
rect 14289 6137 14323 6171
rect 4813 6069 4847 6103
rect 12909 6069 12943 6103
rect 3157 5865 3191 5899
rect 4353 5865 4387 5899
rect 5365 5865 5399 5899
rect 8953 5865 8987 5899
rect 10793 5865 10827 5899
rect 12817 5865 12851 5899
rect 4813 5797 4847 5831
rect 8125 5797 8159 5831
rect 11253 5797 11287 5831
rect 13369 5797 13403 5831
rect 7297 5729 7331 5763
rect 7941 5729 7975 5763
rect 8033 5729 8067 5763
rect 9597 5729 9631 5763
rect 10241 5729 10275 5763
rect 11621 5729 11655 5763
rect 15025 5729 15059 5763
rect 1593 5661 1627 5695
rect 2053 5661 2087 5695
rect 2237 5661 2271 5695
rect 2881 5661 2915 5695
rect 2973 5661 3007 5695
rect 3249 5661 3283 5695
rect 4537 5661 4571 5695
rect 4689 5661 4723 5695
rect 4905 5661 4939 5695
rect 5549 5661 5583 5695
rect 5825 5661 5859 5695
rect 6653 5661 6687 5695
rect 6837 5661 6871 5695
rect 6929 5661 6963 5695
rect 7757 5661 7791 5695
rect 8217 5661 8251 5695
rect 9137 5661 9171 5695
rect 9229 5661 9263 5695
rect 10517 5661 10551 5695
rect 11437 5661 11471 5695
rect 11529 5661 11563 5695
rect 11713 5661 11747 5695
rect 14473 5661 14507 5695
rect 14933 5661 14967 5695
rect 15209 5661 15243 5695
rect 15301 5661 15335 5695
rect 7021 5593 7055 5627
rect 7159 5593 7193 5627
rect 9505 5593 9539 5627
rect 13093 5593 13127 5627
rect 14289 5593 14323 5627
rect 1501 5525 1535 5559
rect 2145 5525 2179 5559
rect 2697 5525 2731 5559
rect 5733 5525 5767 5559
rect 8401 5525 8435 5559
rect 10425 5525 10459 5559
rect 10609 5525 10643 5559
rect 13001 5525 13035 5559
rect 13185 5525 13219 5559
rect 14105 5525 14139 5559
rect 15485 5525 15519 5559
rect 3893 5321 3927 5355
rect 10425 5321 10459 5355
rect 10517 5321 10551 5355
rect 12909 5321 12943 5355
rect 14197 5321 14231 5355
rect 14473 5321 14507 5355
rect 3249 5253 3283 5287
rect 4537 5253 4571 5287
rect 5365 5253 5399 5287
rect 10241 5253 10275 5287
rect 12817 5253 12851 5287
rect 13921 5253 13955 5287
rect 1685 5185 1719 5219
rect 2329 5185 2363 5219
rect 3433 5185 3467 5219
rect 4077 5185 4111 5219
rect 4169 5185 4203 5219
rect 5181 5185 5215 5219
rect 5273 5185 5307 5219
rect 5549 5185 5583 5219
rect 6929 5185 6963 5219
rect 7205 5185 7239 5219
rect 7389 5185 7423 5219
rect 7849 5185 7883 5219
rect 8953 5185 8987 5219
rect 10609 5185 10643 5219
rect 11805 5185 11839 5219
rect 11897 5185 11931 5219
rect 12173 5185 12207 5219
rect 13093 5185 13127 5219
rect 13185 5185 13219 5219
rect 13461 5185 13495 5219
rect 14105 5185 14139 5219
rect 14289 5185 14323 5219
rect 4445 5117 4479 5151
rect 7113 5117 7147 5151
rect 8677 5117 8711 5151
rect 12081 5117 12115 5151
rect 12817 5117 12851 5151
rect 13369 5117 13403 5151
rect 14933 5117 14967 5151
rect 15209 5117 15243 5151
rect 16681 5117 16715 5151
rect 4997 5049 5031 5083
rect 7021 5049 7055 5083
rect 1593 4981 1627 5015
rect 2237 4981 2271 5015
rect 3065 4981 3099 5015
rect 6745 4981 6779 5015
rect 8033 4981 8067 5015
rect 10793 4981 10827 5015
rect 11621 4981 11655 5015
rect 1777 4777 1811 4811
rect 3157 4777 3191 4811
rect 5273 4777 5307 4811
rect 7297 4777 7331 4811
rect 8401 4777 8435 4811
rect 10425 4777 10459 4811
rect 11713 4777 11747 4811
rect 13185 4777 13219 4811
rect 13369 4777 13403 4811
rect 14105 4777 14139 4811
rect 3801 4641 3835 4675
rect 11253 4641 11287 4675
rect 13461 4641 13495 4675
rect 14841 4641 14875 4675
rect 1685 4573 1719 4607
rect 1961 4573 1995 4607
rect 2053 4573 2087 4607
rect 3249 4573 3283 4607
rect 3985 4573 4019 4607
rect 4353 4573 4387 4607
rect 4997 4573 5031 4607
rect 5089 4573 5123 4607
rect 5365 4573 5399 4607
rect 5825 4573 5859 4607
rect 6193 4573 6227 4607
rect 7205 4573 7239 4607
rect 8217 4573 8251 4607
rect 8401 4573 8435 4607
rect 8953 4573 8987 4607
rect 9229 4573 9263 4607
rect 10609 4573 10643 4607
rect 11437 4573 11471 4607
rect 11529 4573 11563 4607
rect 11805 4573 11839 4607
rect 12357 4573 12391 4607
rect 13553 4573 13587 4607
rect 14289 4573 14323 4607
rect 15117 4573 15151 4607
rect 4813 4505 4847 4539
rect 6009 4505 6043 4539
rect 10793 4505 10827 4539
rect 12541 4505 12575 4539
rect 2237 4437 2271 4471
rect 3985 4437 4019 4471
rect 4905 4233 4939 4267
rect 8861 4233 8895 4267
rect 12541 4233 12575 4267
rect 15393 4233 15427 4267
rect 5457 4165 5491 4199
rect 10333 4165 10367 4199
rect 14381 4165 14415 4199
rect 14565 4165 14599 4199
rect 15025 4165 15059 4199
rect 15209 4165 15243 4199
rect 1685 4097 1719 4131
rect 2881 4097 2915 4131
rect 3709 4097 3743 4131
rect 4169 4097 4203 4131
rect 4997 4097 5031 4131
rect 5641 4097 5675 4131
rect 5733 4097 5767 4131
rect 6929 4097 6963 4131
rect 7113 4097 7147 4131
rect 7573 4097 7607 4131
rect 9137 4097 9171 4131
rect 10057 4097 10091 4131
rect 10793 4097 10827 4131
rect 11713 4097 11747 4131
rect 11989 4097 12023 4131
rect 12633 4097 12667 4131
rect 13185 4097 13219 4131
rect 13277 4097 13311 4131
rect 1777 4029 1811 4063
rect 1961 4029 1995 4063
rect 2973 4029 3007 4063
rect 7849 4029 7883 4063
rect 9045 4029 9079 4063
rect 9230 4029 9264 4063
rect 9321 4029 9355 4063
rect 10241 4029 10275 4063
rect 11805 4029 11839 4063
rect 3617 3961 3651 3995
rect 7113 3961 7147 3995
rect 1869 3893 1903 3927
rect 4353 3893 4387 3927
rect 5457 3893 5491 3927
rect 9873 3893 9907 3927
rect 10333 3893 10367 3927
rect 10885 3893 10919 3927
rect 11529 3893 11563 3927
rect 11989 3893 12023 3927
rect 14197 3893 14231 3927
rect 5181 3689 5215 3723
rect 7665 3689 7699 3723
rect 9505 3689 9539 3723
rect 10609 3689 10643 3723
rect 11161 3689 11195 3723
rect 15301 3689 15335 3723
rect 3801 3621 3835 3655
rect 11621 3621 11655 3655
rect 12909 3621 12943 3655
rect 13369 3621 13403 3655
rect 2053 3553 2087 3587
rect 2421 3553 2455 3587
rect 2881 3553 2915 3587
rect 4445 3553 4479 3587
rect 8125 3553 8159 3587
rect 8309 3553 8343 3587
rect 9045 3553 9079 3587
rect 14749 3553 14783 3587
rect 1593 3485 1627 3519
rect 2237 3485 2271 3519
rect 3926 3485 3960 3519
rect 4353 3485 4387 3519
rect 4997 3485 5031 3519
rect 5181 3485 5215 3519
rect 5641 3485 5675 3519
rect 5917 3485 5951 3519
rect 6009 3485 6043 3519
rect 7021 3485 7055 3519
rect 8953 3485 8987 3519
rect 9229 3485 9263 3519
rect 9321 3485 9355 3519
rect 10701 3485 10735 3519
rect 11345 3485 11379 3519
rect 11437 3485 11471 3519
rect 11713 3485 11747 3519
rect 12449 3485 12483 3519
rect 13093 3485 13127 3519
rect 13185 3485 13219 3519
rect 13461 3485 13495 3519
rect 14289 3485 14323 3519
rect 14591 3485 14625 3519
rect 15209 3485 15243 3519
rect 1501 3417 1535 3451
rect 5825 3417 5859 3451
rect 6837 3417 6871 3451
rect 14381 3417 14415 3451
rect 14473 3417 14507 3451
rect 2881 3349 2915 3383
rect 3985 3349 4019 3383
rect 6193 3349 6227 3383
rect 6653 3349 6687 3383
rect 8033 3349 8067 3383
rect 10241 3349 10275 3383
rect 12357 3349 12391 3383
rect 14105 3349 14139 3383
rect 2605 3145 2639 3179
rect 11713 3145 11747 3179
rect 1409 3077 1443 3111
rect 3341 3077 3375 3111
rect 4353 3077 4387 3111
rect 13921 3077 13955 3111
rect 14013 3077 14047 3111
rect 14841 3077 14875 3111
rect 1501 3009 1535 3043
rect 1777 3009 1811 3043
rect 1869 3009 1903 3043
rect 2697 3007 2731 3041
rect 3157 3009 3191 3043
rect 3433 3009 3467 3043
rect 4077 3009 4111 3043
rect 5457 3009 5491 3043
rect 5733 3009 5767 3043
rect 7205 3009 7239 3043
rect 7481 3009 7515 3043
rect 8217 3009 8251 3043
rect 8401 3009 8435 3043
rect 8493 3009 8527 3043
rect 8677 3009 8711 3043
rect 9689 3009 9723 3043
rect 10149 3009 10183 3043
rect 10517 3009 10551 3043
rect 11529 3009 11563 3043
rect 12265 3009 12299 3043
rect 13645 3009 13679 3043
rect 14473 3009 14507 3043
rect 14657 3009 14691 3043
rect 15577 3009 15611 3043
rect 3893 2941 3927 2975
rect 4445 2941 4479 2975
rect 5365 2941 5399 2975
rect 5825 2941 5859 2975
rect 7113 2941 7147 2975
rect 7573 2941 7607 2975
rect 9873 2941 9907 2975
rect 10425 2941 10459 2975
rect 12817 2941 12851 2975
rect 13553 2941 13587 2975
rect 2053 2873 2087 2907
rect 4169 2873 4203 2907
rect 8309 2873 8343 2907
rect 10333 2873 10367 2907
rect 15761 2873 15795 2907
rect 3157 2805 3191 2839
rect 5181 2805 5215 2839
rect 6929 2805 6963 2839
rect 8033 2805 8067 2839
rect 13369 2805 13403 2839
rect 4905 2601 4939 2635
rect 6469 2601 6503 2635
rect 7481 2601 7515 2635
rect 8217 2601 8251 2635
rect 8953 2601 8987 2635
rect 9781 2601 9815 2635
rect 12633 2601 12667 2635
rect 13277 2601 13311 2635
rect 13921 2601 13955 2635
rect 14197 2601 14231 2635
rect 8401 2533 8435 2567
rect 10333 2465 10367 2499
rect 14933 2465 14967 2499
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 2881 2397 2915 2431
rect 4353 2397 4387 2431
rect 4905 2397 4939 2431
rect 5089 2397 5123 2431
rect 5733 2397 5767 2431
rect 6377 2397 6411 2431
rect 6653 2397 6687 2431
rect 6745 2397 6779 2431
rect 7573 2397 7607 2431
rect 8033 2397 8067 2431
rect 8217 2397 8251 2431
rect 9137 2397 9171 2431
rect 9965 2397 9999 2431
rect 10057 2397 10091 2431
rect 12081 2397 12115 2431
rect 12817 2397 12851 2431
rect 13461 2397 13495 2431
rect 13921 2397 13955 2431
rect 14381 2397 14415 2431
rect 14841 2397 14875 2431
rect 2697 2329 2731 2363
rect 4169 2329 4203 2363
rect 9321 2329 9355 2363
rect 10425 2329 10459 2363
rect 15485 2329 15519 2363
rect 15669 2329 15703 2363
rect 5641 2261 5675 2295
rect 6929 2261 6963 2295
rect 11989 2261 12023 2295
<< metal1 >>
rect 1104 17434 16468 17456
rect 1104 17382 6103 17434
rect 6155 17382 6167 17434
rect 6219 17382 6231 17434
rect 6283 17382 6295 17434
rect 6347 17382 11224 17434
rect 11276 17382 11288 17434
rect 11340 17382 11352 17434
rect 11404 17382 11416 17434
rect 11468 17382 16468 17434
rect 1104 17360 16468 17382
rect 14 17280 20 17332
rect 72 17320 78 17332
rect 2593 17323 2651 17329
rect 2593 17320 2605 17323
rect 72 17292 2605 17320
rect 72 17280 78 17292
rect 2593 17289 2605 17292
rect 2639 17289 2651 17323
rect 2593 17283 2651 17289
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 12621 17323 12679 17329
rect 12621 17320 12633 17323
rect 9824 17292 12633 17320
rect 9824 17280 9830 17292
rect 12621 17289 12633 17292
rect 12667 17289 12679 17323
rect 12621 17283 12679 17289
rect 1854 17252 1860 17264
rect 1815 17224 1860 17252
rect 1854 17212 1860 17224
rect 1912 17212 1918 17264
rect 4154 17252 4160 17264
rect 4115 17224 4160 17252
rect 4154 17212 4160 17224
rect 4212 17212 4218 17264
rect 7926 17212 7932 17264
rect 7984 17252 7990 17264
rect 8021 17255 8079 17261
rect 8021 17252 8033 17255
rect 7984 17224 8033 17252
rect 7984 17212 7990 17224
rect 8021 17221 8033 17224
rect 8067 17221 8079 17255
rect 8021 17215 8079 17221
rect 8294 17212 8300 17264
rect 8352 17252 8358 17264
rect 9953 17255 10011 17261
rect 9953 17252 9965 17255
rect 8352 17224 9965 17252
rect 8352 17212 8358 17224
rect 9953 17221 9965 17224
rect 9999 17252 10011 17255
rect 10873 17255 10931 17261
rect 10873 17252 10885 17255
rect 9999 17224 10885 17252
rect 9999 17221 10011 17224
rect 9953 17215 10011 17221
rect 10873 17221 10885 17224
rect 10919 17221 10931 17255
rect 10873 17215 10931 17221
rect 11882 17212 11888 17264
rect 11940 17252 11946 17264
rect 17494 17252 17500 17264
rect 11940 17224 13492 17252
rect 11940 17212 11946 17224
rect 1670 17144 1676 17196
rect 1728 17184 1734 17196
rect 2685 17187 2743 17193
rect 2685 17184 2697 17187
rect 1728 17156 2697 17184
rect 1728 17144 1734 17156
rect 2685 17153 2697 17156
rect 2731 17153 2743 17187
rect 2685 17147 2743 17153
rect 4246 17144 4252 17196
rect 4304 17184 4310 17196
rect 4341 17187 4399 17193
rect 4341 17184 4353 17187
rect 4304 17156 4353 17184
rect 4304 17144 4310 17156
rect 4341 17153 4353 17156
rect 4387 17153 4399 17187
rect 5074 17184 5080 17196
rect 5035 17156 5080 17184
rect 4341 17147 4399 17153
rect 5074 17144 5080 17156
rect 5132 17144 5138 17196
rect 5442 17144 5448 17196
rect 5500 17184 5506 17196
rect 5629 17187 5687 17193
rect 5629 17184 5641 17187
rect 5500 17156 5641 17184
rect 5500 17144 5506 17156
rect 5629 17153 5641 17156
rect 5675 17153 5687 17187
rect 5629 17147 5687 17153
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 6365 17187 6423 17193
rect 6365 17184 6377 17187
rect 5960 17156 6377 17184
rect 5960 17144 5966 17156
rect 6365 17153 6377 17156
rect 6411 17153 6423 17187
rect 8202 17184 8208 17196
rect 8163 17156 8208 17184
rect 6365 17147 6423 17153
rect 8202 17144 8208 17156
rect 8260 17144 8266 17196
rect 9217 17187 9275 17193
rect 9217 17153 9229 17187
rect 9263 17153 9275 17187
rect 9398 17184 9404 17196
rect 9359 17156 9404 17184
rect 9217 17147 9275 17153
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17116 2099 17119
rect 6641 17119 6699 17125
rect 2087 17088 5212 17116
rect 2087 17085 2099 17088
rect 2041 17079 2099 17085
rect 4890 17048 4896 17060
rect 4851 17020 4896 17048
rect 4890 17008 4896 17020
rect 4948 17008 4954 17060
rect 5184 17048 5212 17088
rect 6641 17085 6653 17119
rect 6687 17116 6699 17119
rect 6914 17116 6920 17128
rect 6687 17088 6920 17116
rect 6687 17085 6699 17088
rect 6641 17079 6699 17085
rect 6914 17076 6920 17088
rect 6972 17076 6978 17128
rect 9232 17116 9260 17147
rect 9398 17144 9404 17156
rect 9456 17144 9462 17196
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17184 10195 17187
rect 10318 17184 10324 17196
rect 10183 17156 10324 17184
rect 10183 17153 10195 17156
rect 10137 17147 10195 17153
rect 10318 17144 10324 17156
rect 10376 17144 10382 17196
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17153 10839 17187
rect 11698 17184 11704 17196
rect 11659 17156 11704 17184
rect 10781 17147 10839 17153
rect 9306 17116 9312 17128
rect 9219 17088 9312 17116
rect 9306 17076 9312 17088
rect 9364 17116 9370 17128
rect 10796 17116 10824 17147
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 11790 17144 11796 17196
rect 11848 17184 11854 17196
rect 12066 17184 12072 17196
rect 11848 17156 11893 17184
rect 12027 17156 12072 17184
rect 11848 17144 11854 17156
rect 12066 17144 12072 17156
rect 12124 17144 12130 17196
rect 12158 17144 12164 17196
rect 12216 17184 12222 17196
rect 13464 17193 13492 17224
rect 15028 17224 17500 17252
rect 12713 17187 12771 17193
rect 12713 17184 12725 17187
rect 12216 17156 12725 17184
rect 12216 17144 12222 17156
rect 12713 17153 12725 17156
rect 12759 17153 12771 17187
rect 12713 17147 12771 17153
rect 13449 17187 13507 17193
rect 13449 17153 13461 17187
rect 13495 17153 13507 17187
rect 13449 17147 13507 17153
rect 13814 17144 13820 17196
rect 13872 17184 13878 17196
rect 15028 17193 15056 17224
rect 17494 17212 17500 17224
rect 17552 17212 17558 17264
rect 14277 17187 14335 17193
rect 14277 17184 14289 17187
rect 13872 17156 14289 17184
rect 13872 17144 13878 17156
rect 14277 17153 14289 17156
rect 14323 17153 14335 17187
rect 14277 17147 14335 17153
rect 15013 17187 15071 17193
rect 15013 17153 15025 17187
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 15565 17187 15623 17193
rect 15565 17184 15577 17187
rect 15436 17156 15577 17184
rect 15436 17144 15442 17156
rect 15565 17153 15577 17156
rect 15611 17153 15623 17187
rect 15565 17147 15623 17153
rect 9364 17088 10824 17116
rect 9364 17076 9370 17088
rect 7466 17048 7472 17060
rect 5184 17020 7472 17048
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 12894 17008 12900 17060
rect 12952 17048 12958 17060
rect 14829 17051 14887 17057
rect 14829 17048 14841 17051
rect 12952 17020 14841 17048
rect 12952 17008 12958 17020
rect 14829 17017 14841 17020
rect 14875 17017 14887 17051
rect 15746 17048 15752 17060
rect 15707 17020 15752 17048
rect 14829 17011 14887 17017
rect 15746 17008 15752 17020
rect 15804 17008 15810 17060
rect 5721 16983 5779 16989
rect 5721 16949 5733 16983
rect 5767 16980 5779 16983
rect 6086 16980 6092 16992
rect 5767 16952 6092 16980
rect 5767 16949 5779 16952
rect 5721 16943 5779 16949
rect 6086 16940 6092 16952
rect 6144 16940 6150 16992
rect 8110 16940 8116 16992
rect 8168 16980 8174 16992
rect 9033 16983 9091 16989
rect 9033 16980 9045 16983
rect 8168 16952 9045 16980
rect 8168 16940 8174 16952
rect 9033 16949 9045 16952
rect 9079 16949 9091 16983
rect 9033 16943 9091 16949
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 10321 16983 10379 16989
rect 10321 16980 10333 16983
rect 10284 16952 10333 16980
rect 10284 16940 10290 16952
rect 10321 16949 10333 16952
rect 10367 16949 10379 16983
rect 11514 16980 11520 16992
rect 11475 16952 11520 16980
rect 10321 16943 10379 16949
rect 11514 16940 11520 16952
rect 11572 16940 11578 16992
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 11977 16983 12035 16989
rect 11977 16980 11989 16983
rect 11940 16952 11989 16980
rect 11940 16940 11946 16952
rect 11977 16949 11989 16952
rect 12023 16949 12035 16983
rect 11977 16943 12035 16949
rect 12710 16940 12716 16992
rect 12768 16980 12774 16992
rect 13265 16983 13323 16989
rect 13265 16980 13277 16983
rect 12768 16952 13277 16980
rect 12768 16940 12774 16952
rect 13265 16949 13277 16952
rect 13311 16949 13323 16983
rect 13265 16943 13323 16949
rect 14093 16983 14151 16989
rect 14093 16949 14105 16983
rect 14139 16980 14151 16983
rect 14550 16980 14556 16992
rect 14139 16952 14556 16980
rect 14139 16949 14151 16952
rect 14093 16943 14151 16949
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 1104 16890 16468 16912
rect 1104 16838 3542 16890
rect 3594 16838 3606 16890
rect 3658 16838 3670 16890
rect 3722 16838 3734 16890
rect 3786 16838 8664 16890
rect 8716 16838 8728 16890
rect 8780 16838 8792 16890
rect 8844 16838 8856 16890
rect 8908 16838 13785 16890
rect 13837 16838 13849 16890
rect 13901 16838 13913 16890
rect 13965 16838 13977 16890
rect 14029 16838 16468 16890
rect 1104 16816 16468 16838
rect 2317 16779 2375 16785
rect 2317 16745 2329 16779
rect 2363 16776 2375 16779
rect 5074 16776 5080 16788
rect 2363 16748 5080 16776
rect 2363 16745 2375 16748
rect 2317 16739 2375 16745
rect 5074 16736 5080 16748
rect 5132 16736 5138 16788
rect 8113 16779 8171 16785
rect 8113 16745 8125 16779
rect 8159 16776 8171 16779
rect 8202 16776 8208 16788
rect 8159 16748 8208 16776
rect 8159 16745 8171 16748
rect 8113 16739 8171 16745
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 11790 16736 11796 16788
rect 11848 16776 11854 16788
rect 12161 16779 12219 16785
rect 12161 16776 12173 16779
rect 11848 16748 12173 16776
rect 11848 16736 11854 16748
rect 12161 16745 12173 16748
rect 12207 16745 12219 16779
rect 14645 16779 14703 16785
rect 14645 16776 14657 16779
rect 12161 16739 12219 16745
rect 12544 16748 14657 16776
rect 3050 16668 3056 16720
rect 3108 16708 3114 16720
rect 4065 16711 4123 16717
rect 4065 16708 4077 16711
rect 3108 16680 4077 16708
rect 3108 16668 3114 16680
rect 4065 16677 4077 16680
rect 4111 16677 4123 16711
rect 4801 16711 4859 16717
rect 4801 16708 4813 16711
rect 4065 16671 4123 16677
rect 4356 16680 4813 16708
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16640 2099 16643
rect 2087 16612 2636 16640
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16572 2283 16575
rect 2498 16572 2504 16584
rect 2271 16544 2504 16572
rect 2271 16541 2283 16544
rect 2225 16535 2283 16541
rect 2498 16532 2504 16544
rect 2556 16532 2562 16584
rect 2608 16581 2636 16612
rect 3694 16600 3700 16652
rect 3752 16640 3758 16652
rect 4356 16649 4384 16680
rect 4801 16677 4813 16680
rect 4847 16677 4859 16711
rect 4801 16671 4859 16677
rect 3789 16643 3847 16649
rect 3789 16640 3801 16643
rect 3752 16612 3801 16640
rect 3752 16600 3758 16612
rect 3789 16609 3801 16612
rect 3835 16640 3847 16643
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 3835 16612 4353 16640
rect 3835 16609 3847 16612
rect 3789 16603 3847 16609
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 6273 16643 6331 16649
rect 6273 16609 6285 16643
rect 6319 16640 6331 16643
rect 6917 16643 6975 16649
rect 6917 16640 6929 16643
rect 6319 16612 6929 16640
rect 6319 16609 6331 16612
rect 6273 16603 6331 16609
rect 6917 16609 6929 16612
rect 6963 16640 6975 16643
rect 7098 16640 7104 16652
rect 6963 16612 7104 16640
rect 6963 16609 6975 16612
rect 6917 16603 6975 16609
rect 7098 16600 7104 16612
rect 7156 16640 7162 16652
rect 7377 16643 7435 16649
rect 7377 16640 7389 16643
rect 7156 16612 7389 16640
rect 7156 16600 7162 16612
rect 7377 16609 7389 16612
rect 7423 16609 7435 16643
rect 9033 16643 9091 16649
rect 9033 16640 9045 16643
rect 7377 16603 7435 16609
rect 7576 16612 9045 16640
rect 2593 16575 2651 16581
rect 2593 16541 2605 16575
rect 2639 16574 2651 16575
rect 2639 16572 2673 16574
rect 2774 16572 2780 16584
rect 2639 16544 2780 16572
rect 2639 16541 2651 16544
rect 2593 16535 2651 16541
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 3927 16575 3985 16581
rect 3927 16541 3939 16575
rect 3973 16572 3985 16575
rect 4062 16572 4068 16584
rect 3973 16544 4068 16572
rect 3973 16541 3985 16544
rect 3927 16535 3985 16541
rect 4062 16532 4068 16544
rect 4120 16572 4126 16584
rect 4157 16575 4215 16581
rect 4157 16572 4169 16575
rect 4120 16544 4169 16572
rect 4120 16532 4126 16544
rect 4157 16541 4169 16544
rect 4203 16541 4215 16575
rect 4982 16572 4988 16584
rect 4943 16544 4988 16572
rect 4157 16535 4215 16541
rect 4982 16532 4988 16544
rect 5040 16532 5046 16584
rect 5350 16572 5356 16584
rect 5311 16544 5356 16572
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 5810 16572 5816 16584
rect 5771 16544 5816 16572
rect 5810 16532 5816 16544
rect 5868 16532 5874 16584
rect 6086 16572 6092 16584
rect 6047 16544 6092 16572
rect 6086 16532 6092 16544
rect 6144 16532 6150 16584
rect 7006 16572 7012 16584
rect 6919 16544 7012 16572
rect 7006 16532 7012 16544
rect 7064 16572 7070 16584
rect 7285 16575 7343 16581
rect 7285 16572 7297 16575
rect 7064 16544 7297 16572
rect 7064 16532 7070 16544
rect 7285 16541 7297 16544
rect 7331 16572 7343 16575
rect 7576 16572 7604 16612
rect 9033 16609 9045 16612
rect 9079 16609 9091 16643
rect 9033 16603 9091 16609
rect 9861 16643 9919 16649
rect 9861 16609 9873 16643
rect 9907 16640 9919 16643
rect 10321 16643 10379 16649
rect 10321 16640 10333 16643
rect 9907 16612 10333 16640
rect 9907 16609 9919 16612
rect 9861 16603 9919 16609
rect 10321 16609 10333 16612
rect 10367 16640 10379 16643
rect 10410 16640 10416 16652
rect 10367 16612 10416 16640
rect 10367 16609 10379 16612
rect 10321 16603 10379 16609
rect 7331 16544 7604 16572
rect 8113 16575 8171 16581
rect 7331 16541 7343 16544
rect 7285 16535 7343 16541
rect 8113 16541 8125 16575
rect 8159 16572 8171 16575
rect 8294 16572 8300 16584
rect 8159 16544 8300 16572
rect 8159 16541 8171 16544
rect 8113 16535 8171 16541
rect 8294 16532 8300 16544
rect 8352 16532 8358 16584
rect 8386 16532 8392 16584
rect 8444 16572 8450 16584
rect 9398 16572 9404 16584
rect 8444 16544 8489 16572
rect 9311 16544 9404 16572
rect 8444 16532 8450 16544
rect 9398 16532 9404 16544
rect 9456 16572 9462 16584
rect 9876 16572 9904 16603
rect 10410 16600 10416 16612
rect 10468 16600 10474 16652
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16640 11575 16643
rect 11977 16643 12035 16649
rect 11977 16640 11989 16643
rect 11563 16612 11989 16640
rect 11563 16609 11575 16612
rect 11517 16603 11575 16609
rect 11977 16609 11989 16612
rect 12023 16640 12035 16643
rect 12066 16640 12072 16652
rect 12023 16612 12072 16640
rect 12023 16609 12035 16612
rect 11977 16603 12035 16609
rect 12066 16600 12072 16612
rect 12124 16640 12130 16652
rect 12544 16640 12572 16748
rect 14645 16745 14657 16748
rect 14691 16745 14703 16779
rect 14645 16739 14703 16745
rect 13446 16668 13452 16720
rect 13504 16708 13510 16720
rect 14185 16711 14243 16717
rect 14185 16708 14197 16711
rect 13504 16680 14197 16708
rect 13504 16668 13510 16680
rect 14185 16677 14197 16680
rect 14231 16677 14243 16711
rect 14185 16671 14243 16677
rect 12124 16612 12572 16640
rect 13081 16643 13139 16649
rect 12124 16600 12130 16612
rect 13081 16609 13093 16643
rect 13127 16640 13139 16643
rect 13538 16640 13544 16652
rect 13127 16612 13544 16640
rect 13127 16609 13139 16612
rect 13081 16603 13139 16609
rect 13538 16600 13544 16612
rect 13596 16600 13602 16652
rect 9456 16544 9904 16572
rect 9953 16575 10011 16581
rect 9456 16532 9462 16544
rect 9953 16541 9965 16575
rect 9999 16572 10011 16575
rect 10226 16572 10232 16584
rect 9999 16544 10232 16572
rect 9999 16541 10011 16544
rect 9953 16535 10011 16541
rect 10226 16532 10232 16544
rect 10284 16532 10290 16584
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16572 11667 16575
rect 11882 16572 11888 16584
rect 11655 16544 11888 16572
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 13173 16575 13231 16581
rect 13173 16541 13185 16575
rect 13219 16541 13231 16575
rect 13556 16572 13584 16600
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 13556 16544 14105 16572
rect 13173 16535 13231 16541
rect 14093 16541 14105 16544
rect 14139 16541 14151 16575
rect 14366 16572 14372 16584
rect 14327 16544 14372 16572
rect 14093 16535 14151 16541
rect 2038 16464 2044 16516
rect 2096 16504 2102 16516
rect 4890 16504 4896 16516
rect 2096 16476 4896 16504
rect 2096 16464 2102 16476
rect 4890 16464 4896 16476
rect 4948 16464 4954 16516
rect 5077 16507 5135 16513
rect 5077 16473 5089 16507
rect 5123 16473 5135 16507
rect 5077 16467 5135 16473
rect 5169 16507 5227 16513
rect 5169 16473 5181 16507
rect 5215 16504 5227 16507
rect 6104 16504 6132 16532
rect 9214 16504 9220 16516
rect 5215 16476 6132 16504
rect 7392 16476 8432 16504
rect 9175 16476 9220 16504
rect 5215 16473 5227 16476
rect 5169 16467 5227 16473
rect 2498 16436 2504 16448
rect 2459 16408 2504 16436
rect 2498 16396 2504 16408
rect 2556 16396 2562 16448
rect 5092 16436 5120 16467
rect 5442 16436 5448 16448
rect 5092 16408 5448 16436
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 5626 16396 5632 16448
rect 5684 16436 5690 16448
rect 5905 16439 5963 16445
rect 5905 16436 5917 16439
rect 5684 16408 5917 16436
rect 5684 16396 5690 16408
rect 5905 16405 5917 16408
rect 5951 16436 5963 16439
rect 7392 16436 7420 16476
rect 7558 16436 7564 16448
rect 5951 16408 7420 16436
rect 7519 16408 7564 16436
rect 5951 16405 5963 16408
rect 5905 16399 5963 16405
rect 7558 16396 7564 16408
rect 7616 16396 7622 16448
rect 8294 16436 8300 16448
rect 8255 16408 8300 16436
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 8404 16436 8432 16476
rect 9214 16464 9220 16476
rect 9272 16464 9278 16516
rect 11514 16504 11520 16516
rect 9324 16476 11520 16504
rect 9324 16436 9352 16476
rect 11514 16464 11520 16476
rect 11572 16464 11578 16516
rect 13188 16504 13216 16535
rect 14366 16532 14372 16544
rect 14424 16532 14430 16584
rect 14458 16532 14464 16584
rect 14516 16572 14522 16584
rect 14516 16544 14561 16572
rect 14516 16532 14522 16544
rect 13446 16504 13452 16516
rect 13188 16476 13452 16504
rect 13446 16464 13452 16476
rect 13504 16464 13510 16516
rect 15194 16504 15200 16516
rect 15155 16476 15200 16504
rect 15194 16464 15200 16476
rect 15252 16464 15258 16516
rect 15286 16464 15292 16516
rect 15344 16504 15350 16516
rect 15381 16507 15439 16513
rect 15381 16504 15393 16507
rect 15344 16476 15393 16504
rect 15344 16464 15350 16476
rect 15381 16473 15393 16476
rect 15427 16473 15439 16507
rect 15381 16467 15439 16473
rect 8404 16408 9352 16436
rect 10505 16439 10563 16445
rect 10505 16405 10517 16439
rect 10551 16436 10563 16439
rect 12158 16436 12164 16448
rect 10551 16408 12164 16436
rect 10551 16405 10563 16408
rect 10505 16399 10563 16405
rect 12158 16396 12164 16408
rect 12216 16396 12222 16448
rect 12897 16439 12955 16445
rect 12897 16405 12909 16439
rect 12943 16436 12955 16439
rect 14366 16436 14372 16448
rect 12943 16408 14372 16436
rect 12943 16405 12955 16408
rect 12897 16399 12955 16405
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 15565 16439 15623 16445
rect 15565 16405 15577 16439
rect 15611 16436 15623 16439
rect 15654 16436 15660 16448
rect 15611 16408 15660 16436
rect 15611 16405 15623 16408
rect 15565 16399 15623 16405
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 1104 16346 16468 16368
rect 1104 16294 6103 16346
rect 6155 16294 6167 16346
rect 6219 16294 6231 16346
rect 6283 16294 6295 16346
rect 6347 16294 11224 16346
rect 11276 16294 11288 16346
rect 11340 16294 11352 16346
rect 11404 16294 11416 16346
rect 11468 16294 16468 16346
rect 1104 16272 16468 16294
rect 4893 16235 4951 16241
rect 4893 16201 4905 16235
rect 4939 16232 4951 16235
rect 5350 16232 5356 16244
rect 4939 16204 5356 16232
rect 4939 16201 4951 16204
rect 4893 16195 4951 16201
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 5442 16192 5448 16244
rect 5500 16232 5506 16244
rect 5500 16204 5545 16232
rect 5500 16192 5506 16204
rect 8110 16192 8116 16244
rect 8168 16232 8174 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 8168 16204 8217 16232
rect 8168 16192 8174 16204
rect 8205 16201 8217 16204
rect 8251 16201 8263 16235
rect 8205 16195 8263 16201
rect 9217 16235 9275 16241
rect 9217 16201 9229 16235
rect 9263 16232 9275 16235
rect 9306 16232 9312 16244
rect 9263 16204 9312 16232
rect 9263 16201 9275 16204
rect 9217 16195 9275 16201
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 10410 16192 10416 16244
rect 10468 16232 10474 16244
rect 11517 16235 11575 16241
rect 11517 16232 11529 16235
rect 10468 16204 11529 16232
rect 10468 16192 10474 16204
rect 11517 16201 11529 16204
rect 11563 16201 11575 16235
rect 15378 16232 15384 16244
rect 15339 16204 15384 16232
rect 11517 16195 11575 16201
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 5460 16164 5488 16192
rect 5626 16164 5632 16176
rect 4080 16136 5488 16164
rect 5587 16136 5632 16164
rect 3694 16096 3700 16108
rect 3655 16068 3700 16096
rect 3694 16056 3700 16068
rect 3752 16056 3758 16108
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16096 3847 16099
rect 3970 16096 3976 16108
rect 3835 16068 3976 16096
rect 3835 16065 3847 16068
rect 3789 16059 3847 16065
rect 3970 16056 3976 16068
rect 4028 16056 4034 16108
rect 4080 16105 4108 16136
rect 5626 16124 5632 16136
rect 5684 16124 5690 16176
rect 8128 16164 8156 16192
rect 6840 16136 8156 16164
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16065 4123 16099
rect 4065 16059 4123 16065
rect 4801 16099 4859 16105
rect 4801 16065 4813 16099
rect 4847 16096 4859 16099
rect 4982 16096 4988 16108
rect 4847 16068 4988 16096
rect 4847 16065 4859 16068
rect 4801 16059 4859 16065
rect 4816 16028 4844 16059
rect 4982 16056 4988 16068
rect 5040 16056 5046 16108
rect 5810 16056 5816 16108
rect 5868 16096 5874 16108
rect 6454 16096 6460 16108
rect 5868 16068 6460 16096
rect 5868 16056 5874 16068
rect 6454 16056 6460 16068
rect 6512 16056 6518 16108
rect 6840 16105 6868 16136
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16065 6791 16099
rect 6733 16059 6791 16065
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16065 6883 16099
rect 7098 16096 7104 16108
rect 7059 16068 7104 16096
rect 6825 16059 6883 16065
rect 3988 16000 4844 16028
rect 6748 16028 6776 16059
rect 7098 16056 7104 16068
rect 7156 16056 7162 16108
rect 7929 16099 7987 16105
rect 7929 16065 7941 16099
rect 7975 16096 7987 16099
rect 8128 16096 8156 16136
rect 8294 16124 8300 16176
rect 8352 16164 8358 16176
rect 9401 16167 9459 16173
rect 9401 16164 9413 16167
rect 8352 16136 9413 16164
rect 8352 16124 8358 16136
rect 9401 16133 9413 16136
rect 9447 16164 9459 16167
rect 10137 16167 10195 16173
rect 10137 16164 10149 16167
rect 9447 16136 10149 16164
rect 9447 16133 9459 16136
rect 9401 16127 9459 16133
rect 10137 16133 10149 16136
rect 10183 16133 10195 16167
rect 10137 16127 10195 16133
rect 10505 16167 10563 16173
rect 10505 16133 10517 16167
rect 10551 16164 10563 16167
rect 11054 16164 11060 16176
rect 10551 16136 11060 16164
rect 10551 16133 10563 16136
rect 10505 16127 10563 16133
rect 11054 16124 11060 16136
rect 11112 16124 11118 16176
rect 13541 16167 13599 16173
rect 13541 16133 13553 16167
rect 13587 16164 13599 16167
rect 14366 16164 14372 16176
rect 13587 16136 14372 16164
rect 13587 16133 13599 16136
rect 13541 16127 13599 16133
rect 7975 16068 8156 16096
rect 7975 16065 7987 16068
rect 7929 16059 7987 16065
rect 8386 16056 8392 16108
rect 8444 16096 8450 16108
rect 9585 16099 9643 16105
rect 9585 16096 9597 16099
rect 8444 16068 9597 16096
rect 8444 16056 8450 16068
rect 9585 16065 9597 16068
rect 9631 16096 9643 16099
rect 10318 16096 10324 16108
rect 9631 16068 10180 16096
rect 10279 16068 10324 16096
rect 9631 16065 9643 16068
rect 9585 16059 9643 16065
rect 7558 16028 7564 16040
rect 6748 16000 7564 16028
rect 3988 15904 4016 16000
rect 7558 15988 7564 16000
rect 7616 16028 7622 16040
rect 7745 16031 7803 16037
rect 7745 16028 7757 16031
rect 7616 16000 7757 16028
rect 7616 15988 7622 16000
rect 7745 15997 7757 16000
rect 7791 16028 7803 16031
rect 8297 16031 8355 16037
rect 8297 16028 8309 16031
rect 7791 16000 8309 16028
rect 7791 15997 7803 16000
rect 7745 15991 7803 15997
rect 8297 15997 8309 16000
rect 8343 15997 8355 16031
rect 8297 15991 8355 15997
rect 4062 15920 4068 15972
rect 4120 15960 4126 15972
rect 6549 15963 6607 15969
rect 6549 15960 6561 15963
rect 4120 15932 6561 15960
rect 4120 15920 4126 15932
rect 6549 15929 6561 15932
rect 6595 15929 6607 15963
rect 7006 15960 7012 15972
rect 6967 15932 7012 15960
rect 6549 15923 6607 15929
rect 7006 15920 7012 15932
rect 7064 15920 7070 15972
rect 2498 15852 2504 15904
rect 2556 15892 2562 15904
rect 3513 15895 3571 15901
rect 3513 15892 3525 15895
rect 2556 15864 3525 15892
rect 2556 15852 2562 15864
rect 3513 15861 3525 15864
rect 3559 15861 3571 15895
rect 3970 15892 3976 15904
rect 3931 15864 3976 15892
rect 3513 15855 3571 15861
rect 3970 15852 3976 15864
rect 4028 15852 4034 15904
rect 8021 15895 8079 15901
rect 8021 15861 8033 15895
rect 8067 15892 8079 15895
rect 8202 15892 8208 15904
rect 8067 15864 8208 15892
rect 8067 15861 8079 15864
rect 8021 15855 8079 15861
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 10152 15892 10180 16068
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 10597 16099 10655 16105
rect 10597 16065 10609 16099
rect 10643 16065 10655 16099
rect 11790 16096 11796 16108
rect 11751 16068 11796 16096
rect 10597 16059 10655 16065
rect 10612 15960 10640 16059
rect 11790 16056 11796 16068
rect 11848 16096 11854 16108
rect 12069 16099 12127 16105
rect 12069 16096 12081 16099
rect 11848 16068 12081 16096
rect 11848 16056 11854 16068
rect 12069 16065 12081 16068
rect 12115 16065 12127 16099
rect 12069 16059 12127 16065
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16096 13323 16099
rect 13556 16096 13584 16127
rect 14366 16124 14372 16136
rect 14424 16124 14430 16176
rect 15286 16164 15292 16176
rect 15247 16136 15292 16164
rect 15286 16124 15292 16136
rect 15344 16124 15350 16176
rect 13311 16068 13584 16096
rect 13633 16099 13691 16105
rect 13311 16065 13323 16068
rect 13265 16059 13323 16065
rect 13633 16065 13645 16099
rect 13679 16096 13691 16099
rect 14458 16096 14464 16108
rect 13679 16068 14464 16096
rect 13679 16065 13691 16068
rect 13633 16059 13691 16065
rect 11698 16028 11704 16040
rect 11611 16000 11704 16028
rect 11698 15988 11704 16000
rect 11756 16028 11762 16040
rect 12161 16031 12219 16037
rect 12161 16028 12173 16031
rect 11756 16000 12173 16028
rect 11756 15988 11762 16000
rect 12161 15997 12173 16000
rect 12207 16028 12219 16031
rect 12250 16028 12256 16040
rect 12207 16000 12256 16028
rect 12207 15997 12219 16000
rect 12161 15991 12219 15997
rect 12250 15988 12256 16000
rect 12308 15988 12314 16040
rect 13170 16028 13176 16040
rect 13083 16000 13176 16028
rect 13170 15988 13176 16000
rect 13228 16028 13234 16040
rect 13648 16028 13676 16059
rect 14458 16056 14464 16068
rect 14516 16056 14522 16108
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16065 14611 16099
rect 15194 16096 15200 16108
rect 15155 16068 15200 16096
rect 14553 16059 14611 16065
rect 13228 16000 13676 16028
rect 14568 16028 14596 16059
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 15562 16028 15568 16040
rect 14568 16000 15568 16028
rect 13228 15988 13234 16000
rect 15562 15988 15568 16000
rect 15620 15988 15626 16040
rect 15654 15988 15660 16040
rect 15712 16028 15718 16040
rect 15712 16000 15805 16028
rect 15712 15988 15718 16000
rect 10870 15960 10876 15972
rect 10612 15932 10876 15960
rect 10870 15920 10876 15932
rect 10928 15960 10934 15972
rect 12989 15963 13047 15969
rect 12989 15960 13001 15963
rect 10928 15932 13001 15960
rect 10928 15920 10934 15932
rect 12989 15929 13001 15932
rect 13035 15929 13047 15963
rect 14734 15960 14740 15972
rect 14695 15932 14740 15960
rect 12989 15923 13047 15929
rect 14734 15920 14740 15932
rect 14792 15920 14798 15972
rect 15672 15892 15700 15988
rect 10152 15864 15700 15892
rect 1104 15802 16468 15824
rect 1104 15750 3542 15802
rect 3594 15750 3606 15802
rect 3658 15750 3670 15802
rect 3722 15750 3734 15802
rect 3786 15750 8664 15802
rect 8716 15750 8728 15802
rect 8780 15750 8792 15802
rect 8844 15750 8856 15802
rect 8908 15750 13785 15802
rect 13837 15750 13849 15802
rect 13901 15750 13913 15802
rect 13965 15750 13977 15802
rect 14029 15750 16468 15802
rect 1104 15728 16468 15750
rect 1486 15648 1492 15700
rect 1544 15688 1550 15700
rect 1581 15691 1639 15697
rect 1581 15688 1593 15691
rect 1544 15660 1593 15688
rect 1544 15648 1550 15660
rect 1581 15657 1593 15660
rect 1627 15657 1639 15691
rect 2498 15688 2504 15700
rect 2459 15660 2504 15688
rect 1581 15651 1639 15657
rect 2498 15648 2504 15660
rect 2556 15648 2562 15700
rect 9953 15691 10011 15697
rect 9953 15657 9965 15691
rect 9999 15688 10011 15691
rect 10318 15688 10324 15700
rect 9999 15660 10324 15688
rect 9999 15657 10011 15660
rect 9953 15651 10011 15657
rect 10318 15648 10324 15660
rect 10376 15648 10382 15700
rect 12986 15688 12992 15700
rect 11624 15660 12848 15688
rect 12947 15660 12992 15688
rect 1673 15623 1731 15629
rect 1673 15589 1685 15623
rect 1719 15620 1731 15623
rect 2130 15620 2136 15632
rect 1719 15592 2136 15620
rect 1719 15589 1731 15592
rect 1673 15583 1731 15589
rect 2130 15580 2136 15592
rect 2188 15580 2194 15632
rect 2516 15552 2544 15648
rect 1780 15524 2544 15552
rect 2685 15555 2743 15561
rect 1780 15493 1808 15524
rect 2685 15521 2697 15555
rect 2731 15552 2743 15555
rect 3326 15552 3332 15564
rect 2731 15524 3332 15552
rect 2731 15521 2743 15524
rect 2685 15515 2743 15521
rect 3326 15512 3332 15524
rect 3384 15552 3390 15564
rect 3789 15555 3847 15561
rect 3789 15552 3801 15555
rect 3384 15524 3801 15552
rect 3384 15512 3390 15524
rect 3789 15521 3801 15524
rect 3835 15521 3847 15555
rect 3789 15515 3847 15521
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15453 1823 15487
rect 1765 15447 1823 15453
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15484 2467 15487
rect 2774 15484 2780 15496
rect 2455 15456 2780 15484
rect 2455 15453 2467 15456
rect 2409 15447 2467 15453
rect 1489 15419 1547 15425
rect 1489 15385 1501 15419
rect 1535 15416 1547 15419
rect 2424 15416 2452 15447
rect 2774 15444 2780 15456
rect 2832 15444 2838 15496
rect 9214 15444 9220 15496
rect 9272 15484 9278 15496
rect 9861 15487 9919 15493
rect 9861 15484 9873 15487
rect 9272 15456 9873 15484
rect 9272 15444 9278 15456
rect 9861 15453 9873 15456
rect 9907 15484 9919 15487
rect 10505 15487 10563 15493
rect 10505 15484 10517 15487
rect 9907 15456 10517 15484
rect 9907 15453 9919 15456
rect 9861 15447 9919 15453
rect 10505 15453 10517 15456
rect 10551 15453 10563 15487
rect 10870 15484 10876 15496
rect 10831 15456 10876 15484
rect 10505 15447 10563 15453
rect 10870 15444 10876 15456
rect 10928 15444 10934 15496
rect 11624 15493 11652 15660
rect 12526 15620 12532 15632
rect 12084 15592 12532 15620
rect 12084 15493 12112 15592
rect 12526 15580 12532 15592
rect 12584 15580 12590 15632
rect 12820 15620 12848 15660
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 13170 15688 13176 15700
rect 13131 15660 13176 15688
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 15194 15688 15200 15700
rect 15155 15660 15200 15688
rect 15194 15648 15200 15660
rect 15252 15648 15258 15700
rect 15470 15620 15476 15632
rect 12820 15592 15476 15620
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15453 11667 15487
rect 11609 15447 11667 15453
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15453 12127 15487
rect 12069 15447 12127 15453
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 12713 15487 12771 15493
rect 12713 15484 12725 15487
rect 12308 15456 12725 15484
rect 12308 15444 12314 15456
rect 12713 15453 12725 15456
rect 12759 15453 12771 15487
rect 12713 15447 12771 15453
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15484 14703 15487
rect 14918 15484 14924 15496
rect 14691 15456 14924 15484
rect 14691 15453 14703 15456
rect 14645 15447 14703 15453
rect 14918 15444 14924 15456
rect 14976 15444 14982 15496
rect 15013 15487 15071 15493
rect 15013 15453 15025 15487
rect 15059 15453 15071 15487
rect 15013 15447 15071 15453
rect 1535 15388 2452 15416
rect 1535 15385 1547 15388
rect 1489 15379 1547 15385
rect 3142 15376 3148 15428
rect 3200 15416 3206 15428
rect 3973 15419 4031 15425
rect 3973 15416 3985 15419
rect 3200 15388 3985 15416
rect 3200 15376 3206 15388
rect 3973 15385 3985 15388
rect 4019 15385 4031 15419
rect 4154 15416 4160 15428
rect 4115 15388 4160 15416
rect 3973 15379 4031 15385
rect 4154 15376 4160 15388
rect 4212 15376 4218 15428
rect 10689 15419 10747 15425
rect 10689 15385 10701 15419
rect 10735 15416 10747 15419
rect 11054 15416 11060 15428
rect 10735 15388 11060 15416
rect 10735 15385 10747 15388
rect 10689 15379 10747 15385
rect 11054 15376 11060 15388
rect 11112 15416 11118 15428
rect 12342 15416 12348 15428
rect 11112 15388 12348 15416
rect 11112 15376 11118 15388
rect 12342 15376 12348 15388
rect 12400 15376 12406 15428
rect 14090 15376 14096 15428
rect 14148 15416 14154 15428
rect 14553 15419 14611 15425
rect 14553 15416 14565 15419
rect 14148 15388 14565 15416
rect 14148 15376 14154 15388
rect 14553 15385 14565 15388
rect 14599 15416 14611 15419
rect 15028 15416 15056 15447
rect 14599 15388 15056 15416
rect 14599 15385 14611 15388
rect 14553 15379 14611 15385
rect 2406 15308 2412 15360
rect 2464 15348 2470 15360
rect 2685 15351 2743 15357
rect 2685 15348 2697 15351
rect 2464 15320 2697 15348
rect 2464 15308 2470 15320
rect 2685 15317 2697 15320
rect 2731 15317 2743 15351
rect 2685 15311 2743 15317
rect 10318 15308 10324 15360
rect 10376 15348 10382 15360
rect 11425 15351 11483 15357
rect 11425 15348 11437 15351
rect 10376 15320 11437 15348
rect 10376 15308 10382 15320
rect 11425 15317 11437 15320
rect 11471 15317 11483 15351
rect 11425 15311 11483 15317
rect 12253 15351 12311 15357
rect 12253 15317 12265 15351
rect 12299 15348 12311 15351
rect 14642 15348 14648 15360
rect 12299 15320 14648 15348
rect 12299 15317 12311 15320
rect 12253 15311 12311 15317
rect 14642 15308 14648 15320
rect 14700 15308 14706 15360
rect 1104 15258 16468 15280
rect 1104 15206 6103 15258
rect 6155 15206 6167 15258
rect 6219 15206 6231 15258
rect 6283 15206 6295 15258
rect 6347 15206 11224 15258
rect 11276 15206 11288 15258
rect 11340 15206 11352 15258
rect 11404 15206 11416 15258
rect 11468 15206 16468 15258
rect 1104 15184 16468 15206
rect 3789 15147 3847 15153
rect 3789 15113 3801 15147
rect 3835 15144 3847 15147
rect 3970 15144 3976 15156
rect 3835 15116 3976 15144
rect 3835 15113 3847 15116
rect 3789 15107 3847 15113
rect 3970 15104 3976 15116
rect 4028 15104 4034 15156
rect 6454 15144 6460 15156
rect 6415 15116 6460 15144
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 7837 15147 7895 15153
rect 7837 15113 7849 15147
rect 7883 15113 7895 15147
rect 7837 15107 7895 15113
rect 5537 15079 5595 15085
rect 5537 15076 5549 15079
rect 3988 15048 4476 15076
rect 2133 15011 2191 15017
rect 2133 14977 2145 15011
rect 2179 15008 2191 15011
rect 2406 15008 2412 15020
rect 2179 14980 2412 15008
rect 2179 14977 2191 14980
rect 2133 14971 2191 14977
rect 2406 14968 2412 14980
rect 2464 14968 2470 15020
rect 3326 15008 3332 15020
rect 3287 14980 3332 15008
rect 3326 14968 3332 14980
rect 3384 14968 3390 15020
rect 3988 15017 4016 15048
rect 3973 15011 4031 15017
rect 3973 14977 3985 15011
rect 4019 14977 4031 15011
rect 3973 14971 4031 14977
rect 4065 15011 4123 15017
rect 4065 14977 4077 15011
rect 4111 14977 4123 15011
rect 4065 14971 4123 14977
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14940 2099 14943
rect 2501 14943 2559 14949
rect 2501 14940 2513 14943
rect 2087 14912 2513 14940
rect 2087 14909 2099 14912
rect 2041 14903 2099 14909
rect 2501 14909 2513 14912
rect 2547 14909 2559 14943
rect 4080 14940 4108 14971
rect 4448 14952 4476 15048
rect 5092 15048 5549 15076
rect 4341 14943 4399 14949
rect 4341 14940 4353 14943
rect 4080 14912 4353 14940
rect 2501 14903 2559 14909
rect 4341 14909 4353 14912
rect 4387 14909 4399 14943
rect 4341 14903 4399 14909
rect 2056 14872 2084 14903
rect 2130 14872 2136 14884
rect 2056 14844 2136 14872
rect 2130 14832 2136 14844
rect 2188 14832 2194 14884
rect 4356 14872 4384 14903
rect 4430 14900 4436 14952
rect 4488 14940 4494 14952
rect 4488 14912 4533 14940
rect 4488 14900 4494 14912
rect 4982 14900 4988 14952
rect 5040 14940 5046 14952
rect 5092 14949 5120 15048
rect 5537 15045 5549 15048
rect 5583 15045 5595 15079
rect 7009 15079 7067 15085
rect 7009 15076 7021 15079
rect 5537 15039 5595 15045
rect 6748 15048 7021 15076
rect 6748 15017 6776 15048
rect 7009 15045 7021 15048
rect 7055 15076 7067 15079
rect 7374 15076 7380 15088
rect 7055 15048 7380 15076
rect 7055 15045 7067 15048
rect 7009 15039 7067 15045
rect 7374 15036 7380 15048
rect 7432 15076 7438 15088
rect 7852 15076 7880 15107
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 11940 15116 12173 15144
rect 11940 15104 11946 15116
rect 12161 15113 12173 15116
rect 12207 15113 12219 15147
rect 12161 15107 12219 15113
rect 12342 15104 12348 15156
rect 12400 15144 12406 15156
rect 13633 15147 13691 15153
rect 13633 15144 13645 15147
rect 12400 15116 13645 15144
rect 12400 15104 12406 15116
rect 13633 15113 13645 15116
rect 13679 15113 13691 15147
rect 13633 15107 13691 15113
rect 14918 15104 14924 15156
rect 14976 15144 14982 15156
rect 15289 15147 15347 15153
rect 15289 15144 15301 15147
rect 14976 15116 15301 15144
rect 14976 15104 14982 15116
rect 15289 15113 15301 15116
rect 15335 15113 15347 15147
rect 15289 15107 15347 15113
rect 7432 15048 7880 15076
rect 7432 15036 7438 15048
rect 11606 15036 11612 15088
rect 11664 15076 11670 15088
rect 14936 15076 14964 15104
rect 11664 15048 11928 15076
rect 11664 15036 11670 15048
rect 5169 15011 5227 15017
rect 5169 14977 5181 15011
rect 5215 15008 5227 15011
rect 6733 15011 6791 15017
rect 5215 14980 5488 15008
rect 5215 14977 5227 14980
rect 5169 14971 5227 14977
rect 5460 14952 5488 14980
rect 6733 14977 6745 15011
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 7558 14968 7564 15020
rect 7616 15008 7622 15020
rect 8113 15011 8171 15017
rect 8113 15008 8125 15011
rect 7616 14980 8125 15008
rect 7616 14968 7622 14980
rect 8113 14977 8125 14980
rect 8159 15008 8171 15011
rect 8389 15011 8447 15017
rect 8389 15008 8401 15011
rect 8159 14980 8401 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8389 14977 8401 14980
rect 8435 15008 8447 15011
rect 11330 15008 11336 15020
rect 8435 14980 11336 15008
rect 8435 14977 8447 14980
rect 8389 14971 8447 14977
rect 11330 14968 11336 14980
rect 11388 14968 11394 15020
rect 11900 15017 11928 15048
rect 13924 15048 14964 15076
rect 11517 15011 11575 15017
rect 11517 14977 11529 15011
rect 11563 15008 11575 15011
rect 11885 15011 11943 15017
rect 11563 14980 11836 15008
rect 11563 14977 11575 14980
rect 11517 14971 11575 14977
rect 5077 14943 5135 14949
rect 5077 14940 5089 14943
rect 5040 14912 5089 14940
rect 5040 14900 5046 14912
rect 5077 14909 5089 14912
rect 5123 14909 5135 14943
rect 5442 14940 5448 14952
rect 5403 14912 5448 14940
rect 5077 14903 5135 14909
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14909 6699 14943
rect 6641 14903 6699 14909
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14940 7159 14943
rect 7282 14940 7288 14952
rect 7147 14912 7288 14940
rect 7147 14909 7159 14912
rect 7101 14903 7159 14909
rect 4522 14872 4528 14884
rect 4356 14844 4528 14872
rect 4522 14832 4528 14844
rect 4580 14872 4586 14884
rect 4893 14875 4951 14881
rect 4893 14872 4905 14875
rect 4580 14844 4905 14872
rect 4580 14832 4586 14844
rect 4893 14841 4905 14844
rect 4939 14841 4951 14875
rect 6656 14872 6684 14903
rect 7116 14872 7144 14903
rect 7282 14900 7288 14912
rect 7340 14900 7346 14952
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14909 8079 14943
rect 8021 14903 8079 14909
rect 6656 14844 7144 14872
rect 8036 14872 8064 14903
rect 8478 14900 8484 14952
rect 8536 14940 8542 14952
rect 11606 14940 11612 14952
rect 8536 14912 8581 14940
rect 11567 14912 11612 14940
rect 8536 14900 8542 14912
rect 11606 14900 11612 14912
rect 11664 14900 11670 14952
rect 11808 14940 11836 14980
rect 11885 14977 11897 15011
rect 11931 14977 11943 15011
rect 11885 14971 11943 14977
rect 12621 15011 12679 15017
rect 12621 14977 12633 15011
rect 12667 15008 12679 15011
rect 12710 15008 12716 15020
rect 12667 14980 12716 15008
rect 12667 14977 12679 14980
rect 12621 14971 12679 14977
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 13924 15017 13952 15048
rect 13817 15011 13875 15017
rect 13817 14977 13829 15011
rect 13863 14977 13875 15011
rect 13817 14971 13875 14977
rect 13909 15011 13967 15017
rect 13909 14977 13921 15011
rect 13955 14977 13967 15011
rect 13909 14971 13967 14977
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 15008 14243 15011
rect 14645 15011 14703 15017
rect 14645 15008 14657 15011
rect 14231 14980 14657 15008
rect 14231 14977 14243 14980
rect 14185 14971 14243 14977
rect 14645 14977 14657 14980
rect 14691 15008 14703 15011
rect 15010 15008 15016 15020
rect 14691 14980 14872 15008
rect 14971 14980 15016 15008
rect 14691 14977 14703 14980
rect 14645 14971 14703 14977
rect 11974 14940 11980 14952
rect 11808 14912 11980 14940
rect 11974 14900 11980 14912
rect 12032 14900 12038 14952
rect 13832 14940 13860 14971
rect 14844 14952 14872 14980
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 13998 14940 14004 14952
rect 13832 14912 14004 14940
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 14737 14943 14795 14949
rect 14737 14909 14749 14943
rect 14783 14909 14795 14943
rect 14737 14903 14795 14909
rect 8496 14872 8524 14900
rect 8036 14844 8524 14872
rect 14093 14875 14151 14881
rect 4893 14835 4951 14841
rect 14093 14841 14105 14875
rect 14139 14872 14151 14875
rect 14752 14872 14780 14903
rect 14826 14900 14832 14952
rect 14884 14940 14890 14952
rect 15105 14943 15163 14949
rect 15105 14940 15117 14943
rect 14884 14912 15117 14940
rect 14884 14900 14890 14912
rect 15105 14909 15117 14912
rect 15151 14909 15163 14943
rect 15105 14903 15163 14909
rect 15010 14872 15016 14884
rect 14139 14844 15016 14872
rect 14139 14841 14151 14844
rect 14093 14835 14151 14841
rect 15010 14832 15016 14844
rect 15068 14832 15074 14884
rect 2498 14764 2504 14816
rect 2556 14804 2562 14816
rect 2685 14807 2743 14813
rect 2685 14804 2697 14807
rect 2556 14776 2697 14804
rect 2556 14764 2562 14776
rect 2685 14773 2697 14776
rect 2731 14773 2743 14807
rect 2685 14767 2743 14773
rect 2958 14764 2964 14816
rect 3016 14804 3022 14816
rect 3237 14807 3295 14813
rect 3237 14804 3249 14807
rect 3016 14776 3249 14804
rect 3016 14764 3022 14776
rect 3237 14773 3249 14776
rect 3283 14773 3295 14807
rect 3237 14767 3295 14773
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 12805 14807 12863 14813
rect 12805 14804 12817 14807
rect 12676 14776 12817 14804
rect 12676 14764 12682 14776
rect 12805 14773 12817 14776
rect 12851 14773 12863 14807
rect 12805 14767 12863 14773
rect 1104 14714 16468 14736
rect 1104 14662 3542 14714
rect 3594 14662 3606 14714
rect 3658 14662 3670 14714
rect 3722 14662 3734 14714
rect 3786 14662 8664 14714
rect 8716 14662 8728 14714
rect 8780 14662 8792 14714
rect 8844 14662 8856 14714
rect 8908 14662 13785 14714
rect 13837 14662 13849 14714
rect 13901 14662 13913 14714
rect 13965 14662 13977 14714
rect 14029 14662 16468 14714
rect 1104 14640 16468 14662
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 2832 14572 2877 14600
rect 2832 14560 2838 14572
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 4212 14572 4261 14600
rect 4212 14560 4218 14572
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 4249 14563 4307 14569
rect 4709 14603 4767 14609
rect 4709 14569 4721 14603
rect 4755 14600 4767 14603
rect 5442 14600 5448 14612
rect 4755 14572 5448 14600
rect 4755 14569 4767 14572
rect 4709 14563 4767 14569
rect 5442 14560 5448 14572
rect 5500 14600 5506 14612
rect 7101 14603 7159 14609
rect 7101 14600 7113 14603
rect 5500 14572 7113 14600
rect 5500 14560 5506 14572
rect 7101 14569 7113 14572
rect 7147 14569 7159 14603
rect 7558 14600 7564 14612
rect 7519 14572 7564 14600
rect 7101 14563 7159 14569
rect 7558 14560 7564 14572
rect 7616 14560 7622 14612
rect 8478 14560 8484 14612
rect 8536 14600 8542 14612
rect 8941 14603 8999 14609
rect 8941 14600 8953 14603
rect 8536 14572 8953 14600
rect 8536 14560 8542 14572
rect 8941 14569 8953 14572
rect 8987 14569 8999 14603
rect 11330 14600 11336 14612
rect 11291 14572 11336 14600
rect 8941 14563 8999 14569
rect 11330 14560 11336 14572
rect 11388 14560 11394 14612
rect 11974 14560 11980 14612
rect 12032 14600 12038 14612
rect 12345 14603 12403 14609
rect 12345 14600 12357 14603
rect 12032 14572 12357 14600
rect 12032 14560 12038 14572
rect 12345 14569 12357 14572
rect 12391 14569 12403 14603
rect 14826 14600 14832 14612
rect 14787 14572 14832 14600
rect 12345 14563 12403 14569
rect 14826 14560 14832 14572
rect 14884 14560 14890 14612
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 15381 14603 15439 14609
rect 15381 14600 15393 14603
rect 15344 14572 15393 14600
rect 15344 14560 15350 14572
rect 15381 14569 15393 14572
rect 15427 14569 15439 14603
rect 15381 14563 15439 14569
rect 8496 14464 8524 14560
rect 11992 14532 12020 14560
rect 11532 14504 12020 14532
rect 10962 14464 10968 14476
rect 7668 14436 8524 14464
rect 10704 14436 10968 14464
rect 1946 14396 1952 14408
rect 1907 14368 1952 14396
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2958 14396 2964 14408
rect 2919 14368 2964 14396
rect 2958 14356 2964 14368
rect 3016 14356 3022 14408
rect 3142 14396 3148 14408
rect 3103 14368 3148 14396
rect 3142 14356 3148 14368
rect 3200 14356 3206 14408
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14396 3295 14399
rect 4154 14396 4160 14408
rect 3283 14368 4160 14396
rect 3283 14365 3295 14368
rect 3237 14359 3295 14365
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 4430 14396 4436 14408
rect 4343 14368 4436 14396
rect 4430 14356 4436 14368
rect 4488 14356 4494 14408
rect 4522 14356 4528 14408
rect 4580 14396 4586 14408
rect 4801 14399 4859 14405
rect 4580 14368 4625 14396
rect 4580 14356 4586 14368
rect 4801 14365 4813 14399
rect 4847 14396 4859 14399
rect 4982 14396 4988 14408
rect 4847 14368 4988 14396
rect 4847 14365 4859 14368
rect 4801 14359 4859 14365
rect 4982 14356 4988 14368
rect 5040 14356 5046 14408
rect 7282 14396 7288 14408
rect 7243 14368 7288 14396
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 7668 14405 7696 14436
rect 7653 14399 7711 14405
rect 7432 14368 7477 14396
rect 7432 14356 7438 14368
rect 7653 14365 7665 14399
rect 7699 14365 7711 14399
rect 7653 14359 7711 14365
rect 8018 14356 8024 14408
rect 8076 14396 8082 14408
rect 8113 14399 8171 14405
rect 8113 14396 8125 14399
rect 8076 14368 8125 14396
rect 8076 14356 8082 14368
rect 8113 14365 8125 14368
rect 8159 14365 8171 14399
rect 8294 14396 8300 14408
rect 8255 14368 8300 14396
rect 8113 14359 8171 14365
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 9122 14396 9128 14408
rect 9083 14368 9128 14396
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 9214 14356 9220 14408
rect 9272 14396 9278 14408
rect 10704 14405 10732 14436
rect 10962 14424 10968 14436
rect 11020 14424 11026 14476
rect 11532 14405 11560 14504
rect 11793 14467 11851 14473
rect 11793 14433 11805 14467
rect 11839 14464 11851 14467
rect 11839 14436 12664 14464
rect 11839 14433 11851 14436
rect 11793 14427 11851 14433
rect 9493 14399 9551 14405
rect 9493 14396 9505 14399
rect 9272 14368 9505 14396
rect 9272 14356 9278 14368
rect 9493 14365 9505 14368
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14365 10747 14399
rect 10689 14359 10747 14365
rect 10873 14399 10931 14405
rect 10873 14365 10885 14399
rect 10919 14365 10931 14399
rect 10873 14359 10931 14365
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14365 11575 14399
rect 11517 14359 11575 14365
rect 4448 14328 4476 14356
rect 9140 14328 9168 14356
rect 9585 14331 9643 14337
rect 9585 14328 9597 14331
rect 4448 14300 7236 14328
rect 9140 14300 9597 14328
rect 7208 14272 7236 14300
rect 9585 14297 9597 14300
rect 9631 14297 9643 14331
rect 10888 14328 10916 14359
rect 11606 14356 11612 14408
rect 11664 14396 11670 14408
rect 12636 14405 12664 14436
rect 14182 14424 14188 14476
rect 14240 14464 14246 14476
rect 14277 14467 14335 14473
rect 14277 14464 14289 14467
rect 14240 14436 14289 14464
rect 14240 14424 14246 14436
rect 14277 14433 14289 14436
rect 14323 14433 14335 14467
rect 14277 14427 14335 14433
rect 11885 14399 11943 14405
rect 11664 14368 11709 14396
rect 11664 14356 11670 14368
rect 11885 14365 11897 14399
rect 11931 14396 11943 14399
rect 12529 14399 12587 14405
rect 12529 14396 12541 14399
rect 11931 14368 12541 14396
rect 11931 14365 11943 14368
rect 11885 14359 11943 14365
rect 12529 14365 12541 14368
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 12621 14399 12679 14405
rect 12621 14365 12633 14399
rect 12667 14396 12679 14399
rect 12897 14399 12955 14405
rect 12897 14396 12909 14399
rect 12667 14368 12909 14396
rect 12667 14365 12679 14368
rect 12621 14359 12679 14365
rect 12897 14365 12909 14368
rect 12943 14396 12955 14399
rect 13262 14396 13268 14408
rect 12943 14368 13268 14396
rect 12943 14365 12955 14368
rect 12897 14359 12955 14365
rect 12434 14328 12440 14340
rect 10888 14300 12440 14328
rect 9585 14291 9643 14297
rect 12434 14288 12440 14300
rect 12492 14288 12498 14340
rect 1578 14220 1584 14272
rect 1636 14260 1642 14272
rect 1765 14263 1823 14269
rect 1765 14260 1777 14263
rect 1636 14232 1777 14260
rect 1636 14220 1642 14232
rect 1765 14229 1777 14232
rect 1811 14229 1823 14263
rect 1765 14223 1823 14229
rect 7190 14220 7196 14272
rect 7248 14260 7254 14272
rect 8205 14263 8263 14269
rect 8205 14260 8217 14263
rect 7248 14232 8217 14260
rect 7248 14220 7254 14232
rect 8205 14229 8217 14232
rect 8251 14229 8263 14263
rect 8205 14223 8263 14229
rect 10134 14220 10140 14272
rect 10192 14260 10198 14272
rect 10781 14263 10839 14269
rect 10781 14260 10793 14263
rect 10192 14232 10793 14260
rect 10192 14220 10198 14232
rect 10781 14229 10793 14232
rect 10827 14229 10839 14263
rect 12544 14260 12572 14359
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 14292 14396 14320 14427
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 14292 14368 14565 14396
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 14645 14399 14703 14405
rect 14645 14365 14657 14399
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14396 15623 14399
rect 15654 14396 15660 14408
rect 15611 14368 15660 14396
rect 15611 14365 15623 14368
rect 15565 14359 15623 14365
rect 12989 14331 13047 14337
rect 12989 14297 13001 14331
rect 13035 14297 13047 14331
rect 12989 14291 13047 14297
rect 14185 14331 14243 14337
rect 14185 14297 14197 14331
rect 14231 14328 14243 14331
rect 14366 14328 14372 14340
rect 14231 14300 14372 14328
rect 14231 14297 14243 14300
rect 14185 14291 14243 14297
rect 13004 14260 13032 14291
rect 14366 14288 14372 14300
rect 14424 14328 14430 14340
rect 14660 14328 14688 14359
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 15746 14328 15752 14340
rect 14424 14300 14688 14328
rect 15707 14300 15752 14328
rect 14424 14288 14430 14300
rect 15746 14288 15752 14300
rect 15804 14288 15810 14340
rect 14550 14260 14556 14272
rect 12544 14232 14556 14260
rect 10781 14223 10839 14229
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 1104 14170 16468 14192
rect 1104 14118 6103 14170
rect 6155 14118 6167 14170
rect 6219 14118 6231 14170
rect 6283 14118 6295 14170
rect 6347 14118 11224 14170
rect 11276 14118 11288 14170
rect 11340 14118 11352 14170
rect 11404 14118 11416 14170
rect 11468 14118 16468 14170
rect 1104 14096 16468 14118
rect 2225 14059 2283 14065
rect 2225 14025 2237 14059
rect 2271 14056 2283 14059
rect 2406 14056 2412 14068
rect 2271 14028 2412 14056
rect 2271 14025 2283 14028
rect 2225 14019 2283 14025
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 7193 14059 7251 14065
rect 7193 14025 7205 14059
rect 7239 14056 7251 14059
rect 7282 14056 7288 14068
rect 7239 14028 7288 14056
rect 7239 14025 7251 14028
rect 7193 14019 7251 14025
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 8018 14056 8024 14068
rect 7979 14028 8024 14056
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 10962 14056 10968 14068
rect 8128 14028 10968 14056
rect 1489 13991 1547 13997
rect 1489 13957 1501 13991
rect 1535 13988 1547 13991
rect 5534 13988 5540 14000
rect 1535 13960 5540 13988
rect 1535 13957 1547 13960
rect 1489 13951 1547 13957
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 8036 13988 8064 14016
rect 7392 13960 8064 13988
rect 1578 13920 1584 13932
rect 1539 13892 1584 13920
rect 1578 13880 1584 13892
rect 1636 13880 1642 13932
rect 2222 13923 2280 13929
rect 2222 13889 2234 13923
rect 2268 13920 2280 13923
rect 2685 13923 2743 13929
rect 2268 13892 2636 13920
rect 2268 13889 2280 13892
rect 2222 13883 2280 13889
rect 2608 13852 2636 13892
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 2958 13920 2964 13932
rect 2731 13892 2964 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 3418 13880 3424 13932
rect 3476 13920 3482 13932
rect 3513 13923 3571 13929
rect 3513 13920 3525 13923
rect 3476 13892 3525 13920
rect 3476 13880 3482 13892
rect 3513 13889 3525 13892
rect 3559 13889 3571 13923
rect 3513 13883 3571 13889
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 3786 13920 3792 13932
rect 3651 13892 3792 13920
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 3786 13880 3792 13892
rect 3844 13880 3850 13932
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13920 3939 13923
rect 3970 13920 3976 13932
rect 3927 13892 3976 13920
rect 3927 13889 3939 13892
rect 3881 13883 3939 13889
rect 3970 13880 3976 13892
rect 4028 13880 4034 13932
rect 5074 13920 5080 13932
rect 5035 13892 5080 13920
rect 5074 13880 5080 13892
rect 5132 13880 5138 13932
rect 5169 13923 5227 13929
rect 5169 13889 5181 13923
rect 5215 13920 5227 13923
rect 5258 13920 5264 13932
rect 5215 13892 5264 13920
rect 5215 13889 5227 13892
rect 5169 13883 5227 13889
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 5350 13880 5356 13932
rect 5408 13920 5414 13932
rect 7392 13929 7420 13960
rect 5445 13923 5503 13929
rect 5445 13920 5457 13923
rect 5408 13892 5457 13920
rect 5408 13880 5414 13892
rect 5445 13889 5457 13892
rect 5491 13889 5503 13923
rect 5445 13883 5503 13889
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13889 7435 13923
rect 7377 13883 7435 13889
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13889 7527 13923
rect 7926 13920 7932 13932
rect 7887 13892 7932 13920
rect 7469 13883 7527 13889
rect 3234 13852 3240 13864
rect 2608 13824 3240 13852
rect 3234 13812 3240 13824
rect 3292 13852 3298 13864
rect 3329 13855 3387 13861
rect 3329 13852 3341 13855
rect 3292 13824 3341 13852
rect 3292 13812 3298 13824
rect 3329 13821 3341 13824
rect 3375 13821 3387 13855
rect 7190 13852 7196 13864
rect 7151 13824 7196 13852
rect 3329 13815 3387 13821
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 7484 13852 7512 13883
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 8128 13929 8156 14028
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 11606 14056 11612 14068
rect 11563 14028 11612 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 11606 14016 11612 14028
rect 11664 14016 11670 14068
rect 12894 14056 12900 14068
rect 11808 14028 12900 14056
rect 9953 13991 10011 13997
rect 9953 13988 9965 13991
rect 9508 13960 9965 13988
rect 8113 13923 8171 13929
rect 8113 13889 8125 13923
rect 8159 13889 8171 13923
rect 8113 13883 8171 13889
rect 9508 13864 9536 13960
rect 9953 13957 9965 13960
rect 9999 13957 10011 13991
rect 9953 13951 10011 13957
rect 11808 13932 11836 14028
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 13538 14016 13544 14068
rect 13596 14056 13602 14068
rect 13725 14059 13783 14065
rect 13725 14056 13737 14059
rect 13596 14028 13737 14056
rect 13596 14016 13602 14028
rect 13725 14025 13737 14028
rect 13771 14025 13783 14059
rect 15562 14056 15568 14068
rect 15523 14028 15568 14056
rect 13725 14019 13783 14025
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 11882 13948 11888 14000
rect 11940 13988 11946 14000
rect 11940 13960 11985 13988
rect 11940 13948 11946 13960
rect 12434 13948 12440 14000
rect 12492 13988 12498 14000
rect 13630 13988 13636 14000
rect 12492 13960 13636 13988
rect 12492 13948 12498 13960
rect 13630 13948 13636 13960
rect 13688 13948 13694 14000
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 9861 13923 9919 13929
rect 9861 13920 9873 13923
rect 9640 13892 9873 13920
rect 9640 13880 9646 13892
rect 9861 13889 9873 13892
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13920 11023 13923
rect 11606 13920 11612 13932
rect 11011 13892 11612 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 8294 13852 8300 13864
rect 7484 13824 8300 13852
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 9490 13852 9496 13864
rect 9451 13824 9496 13852
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 10873 13855 10931 13861
rect 10873 13821 10885 13855
rect 10919 13852 10931 13855
rect 11146 13852 11152 13864
rect 10919 13824 11152 13852
rect 10919 13821 10931 13824
rect 10873 13815 10931 13821
rect 11146 13812 11152 13824
rect 11204 13852 11210 13864
rect 11716 13852 11744 13883
rect 11790 13880 11796 13932
rect 11848 13920 11854 13932
rect 11848 13892 11893 13920
rect 11848 13880 11854 13892
rect 11974 13880 11980 13932
rect 12032 13929 12038 13932
rect 12032 13923 12061 13929
rect 12049 13889 12061 13923
rect 12032 13883 12061 13889
rect 12805 13923 12863 13929
rect 12805 13889 12817 13923
rect 12851 13920 12863 13923
rect 12894 13920 12900 13932
rect 12851 13892 12900 13920
rect 12851 13889 12863 13892
rect 12805 13883 12863 13889
rect 12032 13880 12038 13883
rect 12894 13880 12900 13892
rect 12952 13880 12958 13932
rect 13909 13923 13967 13929
rect 13909 13889 13921 13923
rect 13955 13889 13967 13923
rect 14182 13920 14188 13932
rect 14143 13892 14188 13920
rect 13909 13883 13967 13889
rect 11204 13824 11744 13852
rect 12161 13855 12219 13861
rect 11204 13812 11210 13824
rect 12161 13821 12173 13855
rect 12207 13821 12219 13855
rect 13924 13852 13952 13883
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 14366 13920 14372 13932
rect 14327 13892 14372 13920
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 15286 13920 15292 13932
rect 15247 13892 15292 13920
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 15654 13920 15660 13932
rect 15615 13892 15660 13920
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 15746 13880 15752 13932
rect 15804 13920 15810 13932
rect 15804 13892 15849 13920
rect 15804 13880 15810 13892
rect 14274 13852 14280 13864
rect 13924 13824 14280 13852
rect 12161 13815 12219 13821
rect 11606 13744 11612 13796
rect 11664 13784 11670 13796
rect 12176 13784 12204 13815
rect 14274 13812 14280 13824
rect 14332 13812 14338 13864
rect 12342 13784 12348 13796
rect 11664 13756 12348 13784
rect 11664 13744 11670 13756
rect 12342 13744 12348 13756
rect 12400 13744 12406 13796
rect 2038 13716 2044 13728
rect 1999 13688 2044 13716
rect 2038 13676 2044 13688
rect 2096 13676 2102 13728
rect 2590 13716 2596 13728
rect 2551 13688 2596 13716
rect 2590 13676 2596 13688
rect 2648 13676 2654 13728
rect 3789 13719 3847 13725
rect 3789 13685 3801 13719
rect 3835 13716 3847 13719
rect 4062 13716 4068 13728
rect 3835 13688 4068 13716
rect 3835 13685 3847 13688
rect 3789 13679 3847 13685
rect 4062 13676 4068 13688
rect 4120 13716 4126 13728
rect 4893 13719 4951 13725
rect 4893 13716 4905 13719
rect 4120 13688 4905 13716
rect 4120 13676 4126 13688
rect 4893 13685 4905 13688
rect 4939 13685 4951 13719
rect 4893 13679 4951 13685
rect 5166 13676 5172 13728
rect 5224 13716 5230 13728
rect 5353 13719 5411 13725
rect 5353 13716 5365 13719
rect 5224 13688 5365 13716
rect 5224 13676 5230 13688
rect 5353 13685 5365 13688
rect 5399 13685 5411 13719
rect 5353 13679 5411 13685
rect 9214 13676 9220 13728
rect 9272 13716 9278 13728
rect 9309 13719 9367 13725
rect 9309 13716 9321 13719
rect 9272 13688 9321 13716
rect 9272 13676 9278 13688
rect 9309 13685 9321 13688
rect 9355 13685 9367 13719
rect 9309 13679 9367 13685
rect 11330 13676 11336 13728
rect 11388 13716 11394 13728
rect 11882 13716 11888 13728
rect 11388 13688 11888 13716
rect 11388 13676 11394 13688
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 12066 13676 12072 13728
rect 12124 13716 12130 13728
rect 12434 13716 12440 13728
rect 12124 13688 12440 13716
rect 12124 13676 12130 13688
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 12710 13716 12716 13728
rect 12671 13688 12716 13716
rect 12710 13676 12716 13688
rect 12768 13676 12774 13728
rect 1104 13626 16468 13648
rect 1104 13574 3542 13626
rect 3594 13574 3606 13626
rect 3658 13574 3670 13626
rect 3722 13574 3734 13626
rect 3786 13574 8664 13626
rect 8716 13574 8728 13626
rect 8780 13574 8792 13626
rect 8844 13574 8856 13626
rect 8908 13574 13785 13626
rect 13837 13574 13849 13626
rect 13901 13574 13913 13626
rect 13965 13574 13977 13626
rect 14029 13574 16468 13626
rect 1104 13552 16468 13574
rect 2130 13512 2136 13524
rect 2091 13484 2136 13512
rect 2130 13472 2136 13484
rect 2188 13472 2194 13524
rect 2590 13472 2596 13524
rect 2648 13512 2654 13524
rect 3053 13515 3111 13521
rect 3053 13512 3065 13515
rect 2648 13484 3065 13512
rect 2648 13472 2654 13484
rect 3053 13481 3065 13484
rect 3099 13481 3111 13515
rect 3053 13475 3111 13481
rect 3789 13515 3847 13521
rect 3789 13481 3801 13515
rect 3835 13512 3847 13515
rect 3878 13512 3884 13524
rect 3835 13484 3884 13512
rect 3835 13481 3847 13484
rect 3789 13475 3847 13481
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 4982 13512 4988 13524
rect 4943 13484 4988 13512
rect 4982 13472 4988 13484
rect 5040 13472 5046 13524
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 10965 13515 11023 13521
rect 10965 13512 10977 13515
rect 8352 13484 10977 13512
rect 8352 13472 8358 13484
rect 10965 13481 10977 13484
rect 11011 13481 11023 13515
rect 10965 13475 11023 13481
rect 11054 13472 11060 13524
rect 11112 13512 11118 13524
rect 12066 13512 12072 13524
rect 11112 13484 12072 13512
rect 11112 13472 11118 13484
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 12342 13512 12348 13524
rect 12303 13484 12348 13512
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 13541 13515 13599 13521
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 14090 13512 14096 13524
rect 13587 13484 14096 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 14090 13472 14096 13484
rect 14148 13472 14154 13524
rect 14182 13472 14188 13524
rect 14240 13512 14246 13524
rect 14461 13515 14519 13521
rect 14461 13512 14473 13515
rect 14240 13484 14473 13512
rect 14240 13472 14246 13484
rect 14461 13481 14473 13484
rect 14507 13481 14519 13515
rect 14461 13475 14519 13481
rect 2608 13376 2636 13472
rect 9401 13447 9459 13453
rect 9401 13413 9413 13447
rect 9447 13444 9459 13447
rect 9582 13444 9588 13456
rect 9447 13416 9588 13444
rect 9447 13413 9459 13416
rect 9401 13407 9459 13413
rect 9582 13404 9588 13416
rect 9640 13444 9646 13456
rect 14826 13444 14832 13456
rect 9640 13416 14832 13444
rect 9640 13404 9646 13416
rect 14826 13404 14832 13416
rect 14884 13404 14890 13456
rect 11146 13376 11152 13388
rect 2332 13348 2636 13376
rect 11107 13348 11152 13376
rect 2332 13317 2360 13348
rect 11146 13336 11152 13348
rect 11204 13336 11210 13388
rect 11241 13379 11299 13385
rect 11241 13345 11253 13379
rect 11287 13376 11299 13379
rect 11790 13376 11796 13388
rect 11287 13348 11796 13376
rect 11287 13345 11299 13348
rect 11241 13339 11299 13345
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13277 2375 13311
rect 2317 13271 2375 13277
rect 2406 13268 2412 13320
rect 2464 13308 2470 13320
rect 2593 13311 2651 13317
rect 2593 13308 2605 13311
rect 2464 13280 2605 13308
rect 2464 13268 2470 13280
rect 2593 13277 2605 13280
rect 2639 13308 2651 13311
rect 2866 13308 2872 13320
rect 2639 13280 2872 13308
rect 2639 13277 2651 13280
rect 2593 13271 2651 13277
rect 2866 13268 2872 13280
rect 2924 13308 2930 13320
rect 3053 13311 3111 13317
rect 3053 13308 3065 13311
rect 2924 13280 3065 13308
rect 2924 13268 2930 13280
rect 3053 13277 3065 13280
rect 3099 13277 3111 13311
rect 3234 13308 3240 13320
rect 3195 13280 3240 13308
rect 3053 13271 3111 13277
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 3970 13308 3976 13320
rect 3931 13280 3976 13308
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4341 13311 4399 13317
rect 4341 13308 4353 13311
rect 4120 13280 4353 13308
rect 4120 13268 4126 13280
rect 4341 13277 4353 13280
rect 4387 13277 4399 13311
rect 4341 13271 4399 13277
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 5169 13311 5227 13317
rect 5169 13308 5181 13311
rect 5132 13280 5181 13308
rect 5132 13268 5138 13280
rect 5169 13277 5181 13280
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 2501 13243 2559 13249
rect 2501 13209 2513 13243
rect 2547 13240 2559 13243
rect 3252 13240 3280 13268
rect 2547 13212 3280 13240
rect 3988 13240 4016 13268
rect 4433 13243 4491 13249
rect 4433 13240 4445 13243
rect 3988 13212 4445 13240
rect 2547 13209 2559 13212
rect 2501 13203 2559 13209
rect 4433 13209 4445 13212
rect 4479 13209 4491 13243
rect 5184 13240 5212 13271
rect 5258 13268 5264 13320
rect 5316 13308 5322 13320
rect 5537 13311 5595 13317
rect 5537 13308 5549 13311
rect 5316 13280 5549 13308
rect 5316 13268 5322 13280
rect 5537 13277 5549 13280
rect 5583 13277 5595 13311
rect 5537 13271 5595 13277
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13308 7711 13311
rect 8754 13308 8760 13320
rect 7699 13280 8760 13308
rect 7699 13277 7711 13280
rect 7653 13271 7711 13277
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 9122 13308 9128 13320
rect 9083 13280 9128 13308
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 9490 13308 9496 13320
rect 9272 13280 9317 13308
rect 9451 13280 9496 13308
rect 9272 13268 9278 13280
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 10318 13308 10324 13320
rect 10279 13280 10324 13308
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 11330 13308 11336 13320
rect 10888 13280 11336 13308
rect 5442 13240 5448 13252
rect 5184 13212 5448 13240
rect 4433 13203 4491 13209
rect 5442 13200 5448 13212
rect 5500 13240 5506 13252
rect 5629 13243 5687 13249
rect 5629 13240 5641 13243
rect 5500 13212 5641 13240
rect 5500 13200 5506 13212
rect 5629 13209 5641 13212
rect 5675 13209 5687 13243
rect 7834 13240 7840 13252
rect 7795 13212 7840 13240
rect 5629 13203 5687 13209
rect 7834 13200 7840 13212
rect 7892 13200 7898 13252
rect 9398 13200 9404 13252
rect 9456 13240 9462 13252
rect 10888 13240 10916 13280
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 11425 13311 11483 13317
rect 11425 13277 11437 13311
rect 11471 13277 11483 13311
rect 11425 13271 11483 13277
rect 9456 13212 10916 13240
rect 9456 13200 9462 13212
rect 11054 13200 11060 13252
rect 11112 13240 11118 13252
rect 11440 13240 11468 13271
rect 11977 13243 12035 13249
rect 11977 13240 11989 13243
rect 11112 13212 11989 13240
rect 11112 13200 11118 13212
rect 11977 13209 11989 13212
rect 12023 13209 12035 13243
rect 12158 13240 12164 13252
rect 12119 13212 12164 13240
rect 11977 13203 12035 13209
rect 12158 13200 12164 13212
rect 12216 13200 12222 13252
rect 12434 13200 12440 13252
rect 12492 13240 12498 13252
rect 13173 13243 13231 13249
rect 13173 13240 13185 13243
rect 12492 13212 13185 13240
rect 12492 13200 12498 13212
rect 13173 13209 13185 13212
rect 13219 13209 13231 13243
rect 13354 13240 13360 13252
rect 13315 13212 13360 13240
rect 13173 13203 13231 13209
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 7469 13175 7527 13181
rect 7469 13172 7481 13175
rect 7248 13144 7481 13172
rect 7248 13132 7254 13144
rect 7469 13141 7481 13144
rect 7515 13141 7527 13175
rect 8938 13172 8944 13184
rect 8899 13144 8944 13172
rect 7469 13135 7527 13141
rect 8938 13132 8944 13144
rect 8996 13132 9002 13184
rect 10413 13175 10471 13181
rect 10413 13141 10425 13175
rect 10459 13172 10471 13175
rect 10686 13172 10692 13184
rect 10459 13144 10692 13172
rect 10459 13141 10471 13144
rect 10413 13135 10471 13141
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 13188 13172 13216 13203
rect 13354 13200 13360 13212
rect 13412 13200 13418 13252
rect 13538 13200 13544 13252
rect 13596 13240 13602 13252
rect 14093 13243 14151 13249
rect 14093 13240 14105 13243
rect 13596 13212 14105 13240
rect 13596 13200 13602 13212
rect 14093 13209 14105 13212
rect 14139 13209 14151 13243
rect 14274 13240 14280 13252
rect 14235 13212 14280 13240
rect 14093 13203 14151 13209
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 14918 13240 14924 13252
rect 14879 13212 14924 13240
rect 14918 13200 14924 13212
rect 14976 13200 14982 13252
rect 15102 13240 15108 13252
rect 15063 13212 15108 13240
rect 15102 13200 15108 13212
rect 15160 13200 15166 13252
rect 15194 13172 15200 13184
rect 13188 13144 15200 13172
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 15289 13175 15347 13181
rect 15289 13141 15301 13175
rect 15335 13172 15347 13175
rect 15470 13172 15476 13184
rect 15335 13144 15476 13172
rect 15335 13141 15347 13144
rect 15289 13135 15347 13141
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 1104 13082 16468 13104
rect 1104 13030 6103 13082
rect 6155 13030 6167 13082
rect 6219 13030 6231 13082
rect 6283 13030 6295 13082
rect 6347 13030 11224 13082
rect 11276 13030 11288 13082
rect 11340 13030 11352 13082
rect 11404 13030 11416 13082
rect 11468 13030 16468 13082
rect 1104 13008 16468 13030
rect 3142 12928 3148 12980
rect 3200 12968 3206 12980
rect 3421 12971 3479 12977
rect 3421 12968 3433 12971
rect 3200 12940 3433 12968
rect 3200 12928 3206 12940
rect 3421 12937 3433 12940
rect 3467 12937 3479 12971
rect 3421 12931 3479 12937
rect 5169 12971 5227 12977
rect 5169 12937 5181 12971
rect 5215 12968 5227 12971
rect 5258 12968 5264 12980
rect 5215 12940 5264 12968
rect 5215 12937 5227 12940
rect 5169 12931 5227 12937
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 5442 12928 5448 12980
rect 5500 12968 5506 12980
rect 6549 12971 6607 12977
rect 6549 12968 6561 12971
rect 5500 12940 6561 12968
rect 5500 12928 5506 12940
rect 6549 12937 6561 12940
rect 6595 12937 6607 12971
rect 8938 12968 8944 12980
rect 6549 12931 6607 12937
rect 6656 12940 8944 12968
rect 1949 12903 2007 12909
rect 1949 12869 1961 12903
rect 1995 12900 2007 12903
rect 3050 12900 3056 12912
rect 1995 12872 3056 12900
rect 1995 12869 2007 12872
rect 1949 12863 2007 12869
rect 3050 12860 3056 12872
rect 3108 12860 3114 12912
rect 4062 12900 4068 12912
rect 3620 12872 4068 12900
rect 2038 12792 2044 12844
rect 2096 12832 2102 12844
rect 2501 12835 2559 12841
rect 2501 12832 2513 12835
rect 2096 12804 2513 12832
rect 2096 12792 2102 12804
rect 2501 12801 2513 12804
rect 2547 12801 2559 12835
rect 2501 12795 2559 12801
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 1486 12724 1492 12776
rect 1544 12764 1550 12776
rect 2700 12764 2728 12795
rect 3418 12792 3424 12844
rect 3476 12832 3482 12844
rect 3620 12841 3648 12872
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 5721 12903 5779 12909
rect 5721 12900 5733 12903
rect 5460 12872 5733 12900
rect 3605 12835 3663 12841
rect 3605 12832 3617 12835
rect 3476 12804 3617 12832
rect 3476 12792 3482 12804
rect 3605 12801 3617 12804
rect 3651 12801 3663 12835
rect 3605 12795 3663 12801
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 3878 12832 3884 12844
rect 3743 12804 3884 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 3878 12792 3884 12804
rect 3936 12832 3942 12844
rect 3973 12835 4031 12841
rect 3973 12832 3985 12835
rect 3936 12804 3985 12832
rect 3936 12792 3942 12804
rect 3973 12801 3985 12804
rect 4019 12801 4031 12835
rect 3973 12795 4031 12801
rect 5258 12792 5264 12844
rect 5316 12832 5322 12844
rect 5460 12841 5488 12872
rect 5721 12869 5733 12872
rect 5767 12900 5779 12903
rect 6656 12900 6684 12940
rect 8938 12928 8944 12940
rect 8996 12928 9002 12980
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 9401 12971 9459 12977
rect 9401 12968 9413 12971
rect 9180 12940 9413 12968
rect 9180 12928 9186 12940
rect 9401 12937 9413 12940
rect 9447 12937 9459 12971
rect 10870 12968 10876 12980
rect 9401 12931 9459 12937
rect 10060 12940 10876 12968
rect 7190 12900 7196 12912
rect 5767 12872 6684 12900
rect 6748 12872 7196 12900
rect 5767 12869 5779 12872
rect 5721 12863 5779 12869
rect 6748 12841 6776 12872
rect 7190 12860 7196 12872
rect 7248 12860 7254 12912
rect 9306 12860 9312 12912
rect 9364 12900 9370 12912
rect 10060 12900 10088 12940
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 11885 12971 11943 12977
rect 11885 12937 11897 12971
rect 11931 12968 11943 12971
rect 11974 12968 11980 12980
rect 11931 12940 11980 12968
rect 11931 12937 11943 12940
rect 11885 12931 11943 12937
rect 11974 12928 11980 12940
rect 12032 12928 12038 12980
rect 12986 12928 12992 12980
rect 13044 12968 13050 12980
rect 13173 12971 13231 12977
rect 13173 12968 13185 12971
rect 13044 12940 13185 12968
rect 13044 12928 13050 12940
rect 13173 12937 13185 12940
rect 13219 12937 13231 12971
rect 14366 12968 14372 12980
rect 14327 12940 14372 12968
rect 13173 12931 13231 12937
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 15010 12968 15016 12980
rect 14971 12940 15016 12968
rect 15010 12928 15016 12940
rect 15068 12928 15074 12980
rect 10686 12900 10692 12912
rect 9364 12872 10088 12900
rect 10647 12872 10692 12900
rect 9364 12860 9370 12872
rect 10686 12860 10692 12872
rect 10744 12900 10750 12912
rect 11054 12900 11060 12912
rect 10744 12872 11060 12900
rect 10744 12860 10750 12872
rect 11054 12860 11060 12872
rect 11112 12860 11118 12912
rect 14001 12903 14059 12909
rect 14001 12900 14013 12903
rect 11440 12872 14013 12900
rect 11440 12844 11468 12872
rect 14001 12869 14013 12872
rect 14047 12900 14059 12903
rect 14047 12872 14320 12900
rect 14047 12869 14059 12872
rect 14001 12863 14059 12869
rect 5445 12835 5503 12841
rect 5445 12832 5457 12835
rect 5316 12804 5457 12832
rect 5316 12792 5322 12804
rect 5445 12801 5457 12804
rect 5491 12801 5503 12835
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5445 12795 5503 12801
rect 5552 12804 5825 12832
rect 1544 12736 2728 12764
rect 1544 12724 1550 12736
rect 5166 12724 5172 12776
rect 5224 12764 5230 12776
rect 5350 12764 5356 12776
rect 5224 12736 5356 12764
rect 5224 12724 5230 12736
rect 5350 12724 5356 12736
rect 5408 12764 5414 12776
rect 5552 12764 5580 12804
rect 5813 12801 5825 12804
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 6733 12835 6791 12841
rect 6733 12801 6745 12835
rect 6779 12801 6791 12835
rect 6733 12795 6791 12801
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 6871 12804 7144 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 7116 12773 7144 12804
rect 7650 12792 7656 12844
rect 7708 12832 7714 12844
rect 7929 12835 7987 12841
rect 7929 12832 7941 12835
rect 7708 12804 7941 12832
rect 7708 12792 7714 12804
rect 7929 12801 7941 12804
rect 7975 12832 7987 12835
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 7975 12804 8217 12832
rect 7975 12801 7987 12804
rect 7929 12795 7987 12801
rect 8205 12801 8217 12804
rect 8251 12801 8263 12835
rect 8754 12832 8760 12844
rect 8715 12804 8760 12832
rect 8205 12795 8263 12801
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 9674 12832 9680 12844
rect 9635 12804 9680 12832
rect 9674 12792 9680 12804
rect 9732 12832 9738 12844
rect 9953 12835 10011 12841
rect 9953 12832 9965 12835
rect 9732 12804 9965 12832
rect 9732 12792 9738 12804
rect 9953 12801 9965 12804
rect 9999 12801 10011 12835
rect 9953 12795 10011 12801
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 11422 12832 11428 12844
rect 10919 12804 11428 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 11422 12792 11428 12804
rect 11480 12792 11486 12844
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12832 11759 12835
rect 12066 12832 12072 12844
rect 11747 12804 12072 12832
rect 11747 12801 11759 12804
rect 11701 12795 11759 12801
rect 5408 12736 5580 12764
rect 7101 12767 7159 12773
rect 5408 12724 5414 12736
rect 7101 12733 7113 12767
rect 7147 12764 7159 12767
rect 7837 12767 7895 12773
rect 7147 12736 7512 12764
rect 7147 12733 7159 12736
rect 7101 12727 7159 12733
rect 7484 12640 7512 12736
rect 7837 12733 7849 12767
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 7852 12696 7880 12727
rect 8294 12724 8300 12776
rect 8352 12764 8358 12776
rect 8772 12764 8800 12792
rect 9585 12767 9643 12773
rect 8352 12736 8397 12764
rect 8772 12736 9444 12764
rect 8352 12724 8358 12736
rect 8312 12696 8340 12724
rect 7852 12668 8340 12696
rect 9416 12696 9444 12736
rect 9585 12733 9597 12767
rect 9631 12764 9643 12767
rect 9858 12764 9864 12776
rect 9631 12736 9864 12764
rect 9631 12733 9643 12736
rect 9585 12727 9643 12733
rect 9858 12724 9864 12736
rect 9916 12764 9922 12776
rect 10045 12767 10103 12773
rect 10045 12764 10057 12767
rect 9916 12736 10057 12764
rect 9916 12724 9922 12736
rect 10045 12733 10057 12736
rect 10091 12764 10103 12767
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 10091 12736 10517 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 10505 12733 10517 12736
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 11532 12764 11560 12795
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 12434 12792 12440 12844
rect 12492 12832 12498 12844
rect 12621 12835 12679 12841
rect 12621 12832 12633 12835
rect 12492 12804 12633 12832
rect 12492 12792 12498 12804
rect 12621 12801 12633 12804
rect 12667 12801 12679 12835
rect 12894 12832 12900 12844
rect 12855 12804 12900 12832
rect 12621 12795 12679 12801
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12832 13047 12835
rect 13354 12832 13360 12844
rect 13035 12804 13360 12832
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 13354 12792 13360 12804
rect 13412 12792 13418 12844
rect 14182 12832 14188 12844
rect 14143 12804 14188 12832
rect 14182 12792 14188 12804
rect 14240 12792 14246 12844
rect 14292 12832 14320 12872
rect 14366 12832 14372 12844
rect 14292 12804 14372 12832
rect 14366 12792 14372 12804
rect 14424 12792 14430 12844
rect 15102 12792 15108 12844
rect 15160 12832 15166 12844
rect 15197 12835 15255 12841
rect 15197 12832 15209 12835
rect 15160 12804 15209 12832
rect 15160 12792 15166 12804
rect 15197 12801 15209 12804
rect 15243 12801 15255 12835
rect 15470 12832 15476 12844
rect 15431 12804 15476 12832
rect 15197 12795 15255 12801
rect 15212 12764 15240 12795
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 15620 12804 15669 12832
rect 15620 12792 15626 12804
rect 15657 12801 15669 12804
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 16577 12767 16635 12773
rect 16577 12764 16589 12767
rect 11532 12736 12664 12764
rect 15212 12736 16589 12764
rect 11532 12696 11560 12736
rect 12636 12708 12664 12736
rect 16577 12733 16589 12736
rect 16623 12733 16635 12767
rect 16577 12727 16635 12733
rect 9416 12668 11560 12696
rect 12618 12656 12624 12708
rect 12676 12696 12682 12708
rect 12713 12699 12771 12705
rect 12713 12696 12725 12699
rect 12676 12668 12725 12696
rect 12676 12656 12682 12668
rect 12713 12665 12725 12668
rect 12759 12696 12771 12699
rect 13170 12696 13176 12708
rect 12759 12668 13176 12696
rect 12759 12665 12771 12668
rect 12713 12659 12771 12665
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 1854 12628 1860 12640
rect 1815 12600 1860 12628
rect 1854 12588 1860 12600
rect 1912 12588 1918 12640
rect 2038 12588 2044 12640
rect 2096 12628 2102 12640
rect 2501 12631 2559 12637
rect 2501 12628 2513 12631
rect 2096 12600 2513 12628
rect 2096 12588 2102 12600
rect 2501 12597 2513 12600
rect 2547 12597 2559 12631
rect 2501 12591 2559 12597
rect 7466 12588 7472 12640
rect 7524 12628 7530 12640
rect 7653 12631 7711 12637
rect 7653 12628 7665 12631
rect 7524 12600 7665 12628
rect 7524 12588 7530 12600
rect 7653 12597 7665 12600
rect 7699 12597 7711 12631
rect 7653 12591 7711 12597
rect 8941 12631 8999 12637
rect 8941 12597 8953 12631
rect 8987 12628 8999 12631
rect 9306 12628 9312 12640
rect 8987 12600 9312 12628
rect 8987 12597 8999 12600
rect 8941 12591 8999 12597
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 9490 12588 9496 12640
rect 9548 12628 9554 12640
rect 15010 12628 15016 12640
rect 9548 12600 15016 12628
rect 9548 12588 9554 12600
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 1104 12538 16468 12560
rect 1104 12486 3542 12538
rect 3594 12486 3606 12538
rect 3658 12486 3670 12538
rect 3722 12486 3734 12538
rect 3786 12486 8664 12538
rect 8716 12486 8728 12538
rect 8780 12486 8792 12538
rect 8844 12486 8856 12538
rect 8908 12486 13785 12538
rect 13837 12486 13849 12538
rect 13901 12486 13913 12538
rect 13965 12486 13977 12538
rect 14029 12486 16468 12538
rect 1104 12464 16468 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 1670 12424 1676 12436
rect 1627 12396 1676 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 1670 12384 1676 12396
rect 1728 12384 1734 12436
rect 1946 12424 1952 12436
rect 1872 12396 1952 12424
rect 1762 12316 1768 12368
rect 1820 12356 1826 12368
rect 1872 12365 1900 12396
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 7193 12427 7251 12433
rect 7193 12424 7205 12427
rect 4120 12396 7205 12424
rect 4120 12384 4126 12396
rect 7193 12393 7205 12396
rect 7239 12393 7251 12427
rect 7193 12387 7251 12393
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 7834 12424 7840 12436
rect 7340 12396 7840 12424
rect 7340 12384 7346 12396
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 11422 12384 11428 12436
rect 11480 12424 11486 12436
rect 11609 12427 11667 12433
rect 11609 12424 11621 12427
rect 11480 12396 11621 12424
rect 11480 12384 11486 12396
rect 11609 12393 11621 12396
rect 11655 12393 11667 12427
rect 12250 12424 12256 12436
rect 12211 12396 12256 12424
rect 11609 12387 11667 12393
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 12710 12424 12716 12436
rect 12671 12396 12716 12424
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 14182 12384 14188 12436
rect 14240 12424 14246 12436
rect 14645 12427 14703 12433
rect 14240 12396 14596 12424
rect 14240 12384 14246 12396
rect 1857 12359 1915 12365
rect 1857 12356 1869 12359
rect 1820 12328 1869 12356
rect 1820 12316 1826 12328
rect 1857 12325 1869 12328
rect 1903 12325 1915 12359
rect 1857 12319 1915 12325
rect 10594 12316 10600 12368
rect 10652 12356 10658 12368
rect 14458 12356 14464 12368
rect 10652 12328 13492 12356
rect 10652 12316 10658 12328
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 2130 12288 2136 12300
rect 1995 12260 2136 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 2130 12248 2136 12260
rect 2188 12288 2194 12300
rect 2777 12291 2835 12297
rect 2777 12288 2789 12291
rect 2188 12260 2789 12288
rect 2188 12248 2194 12260
rect 2777 12257 2789 12260
rect 2823 12257 2835 12291
rect 7650 12288 7656 12300
rect 7611 12260 7656 12288
rect 2777 12251 2835 12257
rect 7650 12248 7656 12260
rect 7708 12248 7714 12300
rect 8294 12288 8300 12300
rect 7760 12260 8300 12288
rect 1486 12180 1492 12232
rect 1544 12220 1550 12232
rect 1765 12223 1823 12229
rect 1765 12220 1777 12223
rect 1544 12192 1777 12220
rect 1544 12180 1550 12192
rect 1765 12189 1777 12192
rect 1811 12189 1823 12223
rect 2038 12220 2044 12232
rect 1999 12192 2044 12220
rect 1765 12183 1823 12189
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 2222 12220 2228 12232
rect 2183 12192 2228 12220
rect 2222 12180 2228 12192
rect 2280 12220 2286 12232
rect 2869 12223 2927 12229
rect 2869 12220 2881 12223
rect 2280 12192 2881 12220
rect 2280 12180 2286 12192
rect 2869 12189 2881 12192
rect 2915 12189 2927 12223
rect 2869 12183 2927 12189
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7377 12223 7435 12229
rect 7377 12220 7389 12223
rect 7248 12192 7389 12220
rect 7248 12180 7254 12192
rect 7377 12189 7389 12192
rect 7423 12189 7435 12223
rect 7377 12183 7435 12189
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 7760 12229 7788 12260
rect 8294 12248 8300 12260
rect 8352 12288 8358 12300
rect 9217 12291 9275 12297
rect 9217 12288 9229 12291
rect 8352 12260 9229 12288
rect 8352 12248 8358 12260
rect 9217 12257 9229 12260
rect 9263 12257 9275 12291
rect 9217 12251 9275 12257
rect 10873 12291 10931 12297
rect 10873 12257 10885 12291
rect 10919 12288 10931 12291
rect 10919 12260 11928 12288
rect 10919 12257 10931 12260
rect 10873 12251 10931 12257
rect 7745 12223 7803 12229
rect 7524 12192 7569 12220
rect 7524 12180 7530 12192
rect 7745 12189 7757 12223
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12189 8263 12223
rect 8205 12183 8263 12189
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12189 9459 12223
rect 9674 12220 9680 12232
rect 9635 12192 9680 12220
rect 9401 12183 9459 12189
rect 5534 12112 5540 12164
rect 5592 12152 5598 12164
rect 5994 12152 6000 12164
rect 5592 12124 6000 12152
rect 5592 12112 5598 12124
rect 5994 12112 6000 12124
rect 6052 12152 6058 12164
rect 8220 12152 8248 12183
rect 6052 12124 8248 12152
rect 9416 12152 9444 12183
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 9858 12220 9864 12232
rect 9819 12192 9864 12220
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 11054 12180 11060 12232
rect 11112 12220 11118 12232
rect 11149 12223 11207 12229
rect 11149 12220 11161 12223
rect 11112 12192 11161 12220
rect 11112 12180 11118 12192
rect 11149 12189 11161 12192
rect 11195 12189 11207 12223
rect 11790 12220 11796 12232
rect 11751 12192 11796 12220
rect 11149 12183 11207 12189
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 11900 12220 11928 12260
rect 11974 12248 11980 12300
rect 12032 12288 12038 12300
rect 12621 12291 12679 12297
rect 12621 12288 12633 12291
rect 12032 12260 12633 12288
rect 12032 12248 12038 12260
rect 12621 12257 12633 12260
rect 12667 12288 12679 12291
rect 13354 12288 13360 12300
rect 12667 12260 13360 12288
rect 12667 12257 12679 12260
rect 12621 12251 12679 12257
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 13464 12288 13492 12328
rect 13740 12328 14464 12356
rect 13740 12288 13768 12328
rect 14458 12316 14464 12328
rect 14516 12316 14522 12368
rect 14568 12356 14596 12396
rect 14645 12393 14657 12427
rect 14691 12424 14703 12427
rect 14918 12424 14924 12436
rect 14691 12396 14924 12424
rect 14691 12393 14703 12396
rect 14645 12387 14703 12393
rect 14918 12384 14924 12396
rect 14976 12384 14982 12436
rect 15654 12384 15660 12436
rect 15712 12424 15718 12436
rect 15749 12427 15807 12433
rect 15749 12424 15761 12427
rect 15712 12396 15761 12424
rect 15712 12384 15718 12396
rect 15749 12393 15761 12396
rect 15795 12393 15807 12427
rect 15749 12387 15807 12393
rect 14568 12328 14688 12356
rect 14660 12300 14688 12328
rect 14182 12288 14188 12300
rect 13464 12260 13768 12288
rect 14143 12260 14188 12288
rect 14182 12248 14188 12260
rect 14240 12248 14246 12300
rect 14642 12248 14648 12300
rect 14700 12248 14706 12300
rect 12066 12220 12072 12232
rect 11900 12192 12072 12220
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 13170 12220 13176 12232
rect 12492 12192 12537 12220
rect 13131 12192 13176 12220
rect 12492 12180 12498 12192
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 13722 12180 13728 12232
rect 13780 12220 13786 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13780 12192 14105 12220
rect 13780 12180 13786 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14366 12220 14372 12232
rect 14327 12192 14372 12220
rect 14093 12183 14151 12189
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 14458 12180 14464 12232
rect 14516 12220 14522 12232
rect 15197 12223 15255 12229
rect 14516 12192 14561 12220
rect 14516 12180 14522 12192
rect 15197 12189 15209 12223
rect 15243 12220 15255 12223
rect 15470 12220 15476 12232
rect 15243 12192 15476 12220
rect 15243 12189 15255 12192
rect 15197 12183 15255 12189
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 15562 12180 15568 12232
rect 15620 12220 15626 12232
rect 15620 12192 15713 12220
rect 15620 12180 15626 12192
rect 9766 12152 9772 12164
rect 9416 12124 9772 12152
rect 6052 12112 6058 12124
rect 9766 12112 9772 12124
rect 9824 12112 9830 12164
rect 11422 12112 11428 12164
rect 11480 12152 11486 12164
rect 12713 12155 12771 12161
rect 12713 12152 12725 12155
rect 11480 12124 12725 12152
rect 11480 12112 11486 12124
rect 12713 12121 12725 12124
rect 12759 12121 12771 12155
rect 12713 12115 12771 12121
rect 13357 12155 13415 12161
rect 13357 12121 13369 12155
rect 13403 12121 13415 12155
rect 13357 12115 13415 12121
rect 13541 12155 13599 12161
rect 13541 12121 13553 12155
rect 13587 12152 13599 12155
rect 15105 12155 15163 12161
rect 15105 12152 15117 12155
rect 13587 12124 15117 12152
rect 13587 12121 13599 12124
rect 13541 12115 13599 12121
rect 15105 12121 15117 12124
rect 15151 12152 15163 12155
rect 15580 12152 15608 12180
rect 15151 12124 15608 12152
rect 15151 12121 15163 12124
rect 15105 12115 15163 12121
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 8386 12084 8392 12096
rect 8076 12056 8392 12084
rect 8076 12044 8082 12056
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 13372 12084 13400 12115
rect 14642 12084 14648 12096
rect 13372 12056 14648 12084
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 1104 11994 16468 12016
rect 1104 11942 6103 11994
rect 6155 11942 6167 11994
rect 6219 11942 6231 11994
rect 6283 11942 6295 11994
rect 6347 11942 11224 11994
rect 11276 11942 11288 11994
rect 11340 11942 11352 11994
rect 11404 11942 11416 11994
rect 11468 11942 16468 11994
rect 1104 11920 16468 11942
rect 2866 11880 2872 11892
rect 2827 11852 2872 11880
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 3970 11880 3976 11892
rect 3931 11852 3976 11880
rect 3970 11840 3976 11852
rect 4028 11840 4034 11892
rect 5166 11880 5172 11892
rect 5127 11852 5172 11880
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 7650 11840 7656 11892
rect 7708 11880 7714 11892
rect 8021 11883 8079 11889
rect 8021 11880 8033 11883
rect 7708 11852 8033 11880
rect 7708 11840 7714 11852
rect 8021 11849 8033 11852
rect 8067 11849 8079 11883
rect 9674 11880 9680 11892
rect 9635 11852 9680 11880
rect 8021 11843 8079 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 12158 11880 12164 11892
rect 12119 11852 12164 11880
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 14277 11883 14335 11889
rect 14277 11880 14289 11883
rect 13596 11852 14289 11880
rect 13596 11840 13602 11852
rect 14277 11849 14289 11852
rect 14323 11849 14335 11883
rect 14277 11843 14335 11849
rect 15657 11883 15715 11889
rect 15657 11849 15669 11883
rect 15703 11880 15715 11883
rect 15746 11880 15752 11892
rect 15703 11852 15752 11880
rect 15703 11849 15715 11852
rect 15657 11843 15715 11849
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 2130 11772 2136 11824
rect 2188 11812 2194 11824
rect 5626 11812 5632 11824
rect 2188 11784 2268 11812
rect 2188 11772 2194 11784
rect 1762 11704 1768 11756
rect 1820 11744 1826 11756
rect 2240 11753 2268 11784
rect 4172 11784 4660 11812
rect 4172 11753 4200 11784
rect 2041 11747 2099 11753
rect 2041 11744 2053 11747
rect 1820 11716 2053 11744
rect 1820 11704 1826 11716
rect 2041 11713 2053 11716
rect 2087 11713 2099 11747
rect 2041 11707 2099 11713
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11713 2283 11747
rect 2225 11707 2283 11713
rect 3145 11747 3203 11753
rect 3145 11713 3157 11747
rect 3191 11744 3203 11747
rect 4157 11747 4215 11753
rect 3191 11716 3464 11744
rect 3191 11713 3203 11716
rect 3145 11707 3203 11713
rect 3436 11688 3464 11716
rect 4157 11713 4169 11747
rect 4203 11713 4215 11747
rect 4157 11707 4215 11713
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 2133 11679 2191 11685
rect 2133 11645 2145 11679
rect 2179 11645 2191 11679
rect 2133 11639 2191 11645
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11676 2375 11679
rect 2958 11676 2964 11688
rect 2363 11648 2964 11676
rect 2363 11645 2375 11648
rect 2317 11639 2375 11645
rect 2148 11608 2176 11639
rect 2958 11636 2964 11648
rect 3016 11636 3022 11688
rect 3053 11679 3111 11685
rect 3053 11645 3065 11679
rect 3099 11645 3111 11679
rect 3418 11676 3424 11688
rect 3379 11648 3424 11676
rect 3053 11639 3111 11645
rect 2774 11608 2780 11620
rect 2148 11580 2780 11608
rect 2774 11568 2780 11580
rect 2832 11568 2838 11620
rect 2866 11568 2872 11620
rect 2924 11608 2930 11620
rect 3068 11608 3096 11639
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 3513 11679 3571 11685
rect 3513 11645 3525 11679
rect 3559 11645 3571 11679
rect 4264 11676 4292 11707
rect 4632 11688 4660 11784
rect 5368 11784 5632 11812
rect 5368 11753 5396 11784
rect 5626 11772 5632 11784
rect 5684 11812 5690 11824
rect 5813 11815 5871 11821
rect 5813 11812 5825 11815
rect 5684 11784 5825 11812
rect 5684 11772 5690 11784
rect 5813 11781 5825 11784
rect 5859 11781 5871 11815
rect 7926 11812 7932 11824
rect 5813 11775 5871 11781
rect 7116 11784 7932 11812
rect 5353 11747 5411 11753
rect 5353 11713 5365 11747
rect 5399 11713 5411 11747
rect 5353 11707 5411 11713
rect 5445 11747 5503 11753
rect 5445 11713 5457 11747
rect 5491 11744 5503 11747
rect 5491 11716 5764 11744
rect 5491 11713 5503 11716
rect 5445 11707 5503 11713
rect 5736 11688 5764 11716
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 7116 11753 7144 11784
rect 7926 11772 7932 11784
rect 7984 11812 7990 11824
rect 7984 11784 8340 11812
rect 7984 11772 7990 11784
rect 7101 11747 7159 11753
rect 7101 11744 7113 11747
rect 6972 11716 7113 11744
rect 6972 11704 6978 11716
rect 7101 11713 7113 11716
rect 7147 11713 7159 11747
rect 7101 11707 7159 11713
rect 7190 11704 7196 11756
rect 7248 11744 7254 11756
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 7248 11716 7297 11744
rect 7248 11704 7254 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 7466 11704 7472 11756
rect 7524 11744 7530 11756
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 7524 11716 7573 11744
rect 7524 11704 7530 11716
rect 7561 11713 7573 11716
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 4522 11676 4528 11688
rect 4264 11648 4528 11676
rect 3513 11639 3571 11645
rect 3528 11608 3556 11639
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 4614 11636 4620 11688
rect 4672 11676 4678 11688
rect 5718 11676 5724 11688
rect 4672 11648 4717 11676
rect 5679 11648 5724 11676
rect 4672 11636 4678 11648
rect 5718 11636 5724 11648
rect 5776 11636 5782 11688
rect 7374 11636 7380 11688
rect 7432 11676 7438 11688
rect 7432 11648 7477 11676
rect 7432 11636 7438 11648
rect 6917 11611 6975 11617
rect 6917 11608 6929 11611
rect 2924 11580 6929 11608
rect 2924 11568 2930 11580
rect 6917 11577 6929 11580
rect 6963 11577 6975 11611
rect 6917 11571 6975 11577
rect 7193 11611 7251 11617
rect 7193 11577 7205 11611
rect 7239 11608 7251 11611
rect 8110 11608 8116 11620
rect 7239 11580 8116 11608
rect 7239 11577 7251 11580
rect 7193 11571 7251 11577
rect 8110 11568 8116 11580
rect 8168 11568 8174 11620
rect 8220 11608 8248 11707
rect 8312 11676 8340 11784
rect 8386 11772 8392 11824
rect 8444 11812 8450 11824
rect 9309 11815 9367 11821
rect 8444 11784 8489 11812
rect 8444 11772 8450 11784
rect 9309 11781 9321 11815
rect 9355 11812 9367 11815
rect 9766 11812 9772 11824
rect 9355 11784 9772 11812
rect 9355 11781 9367 11784
rect 9309 11775 9367 11781
rect 9766 11772 9772 11784
rect 9824 11772 9830 11824
rect 14182 11812 14188 11824
rect 9876 11784 14188 11812
rect 9490 11744 9496 11756
rect 9451 11716 9496 11744
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 9876 11676 9904 11784
rect 14182 11772 14188 11784
rect 14240 11772 14246 11824
rect 15102 11772 15108 11824
rect 15160 11812 15166 11824
rect 15197 11815 15255 11821
rect 15197 11812 15209 11815
rect 15160 11784 15209 11812
rect 15160 11772 15166 11784
rect 15197 11781 15209 11784
rect 15243 11781 15255 11815
rect 15197 11775 15255 11781
rect 10318 11704 10324 11756
rect 10376 11744 10382 11756
rect 10965 11747 11023 11753
rect 10965 11744 10977 11747
rect 10376 11716 10977 11744
rect 10376 11704 10382 11716
rect 10965 11713 10977 11716
rect 11011 11713 11023 11747
rect 11606 11744 11612 11756
rect 11567 11716 11612 11744
rect 10965 11707 11023 11713
rect 11606 11704 11612 11716
rect 11664 11704 11670 11756
rect 11882 11744 11888 11756
rect 11843 11716 11888 11744
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 11974 11704 11980 11756
rect 12032 11744 12038 11756
rect 12805 11747 12863 11753
rect 12032 11716 12077 11744
rect 12032 11704 12038 11716
rect 12805 11713 12817 11747
rect 12851 11744 12863 11747
rect 13078 11744 13084 11756
rect 12851 11716 13084 11744
rect 12851 11713 12863 11716
rect 12805 11707 12863 11713
rect 13078 11704 13084 11716
rect 13136 11704 13142 11756
rect 13722 11744 13728 11756
rect 13635 11716 13728 11744
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 13998 11744 14004 11756
rect 13959 11716 14004 11744
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14093 11747 14151 11753
rect 14093 11713 14105 11747
rect 14139 11713 14151 11747
rect 14093 11707 14151 11713
rect 10686 11676 10692 11688
rect 8312 11648 9904 11676
rect 10647 11648 10692 11676
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 11701 11679 11759 11685
rect 11701 11645 11713 11679
rect 11747 11676 11759 11679
rect 11790 11676 11796 11688
rect 11747 11648 11796 11676
rect 11747 11645 11759 11648
rect 11701 11639 11759 11645
rect 11790 11636 11796 11648
rect 11848 11676 11854 11688
rect 12713 11679 12771 11685
rect 12713 11676 12725 11679
rect 11848 11648 12725 11676
rect 11848 11636 11854 11648
rect 12713 11645 12725 11648
rect 12759 11645 12771 11679
rect 13740 11676 13768 11704
rect 14108 11676 14136 11707
rect 14918 11704 14924 11756
rect 14976 11744 14982 11756
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 14976 11716 15485 11744
rect 14976 11704 14982 11716
rect 15473 11713 15485 11716
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 14458 11676 14464 11688
rect 13740 11648 13952 11676
rect 14108 11648 14464 11676
rect 12713 11639 12771 11645
rect 8478 11608 8484 11620
rect 8220 11580 8484 11608
rect 8478 11568 8484 11580
rect 8536 11608 8542 11620
rect 12066 11608 12072 11620
rect 8536 11580 12072 11608
rect 8536 11568 8542 11580
rect 12066 11568 12072 11580
rect 12124 11568 12130 11620
rect 13354 11568 13360 11620
rect 13412 11608 13418 11620
rect 13817 11611 13875 11617
rect 13817 11608 13829 11611
rect 13412 11580 13829 11608
rect 13412 11568 13418 11580
rect 13817 11577 13829 11580
rect 13863 11577 13875 11611
rect 13817 11571 13875 11577
rect 1857 11543 1915 11549
rect 1857 11509 1869 11543
rect 1903 11540 1915 11543
rect 2130 11540 2136 11552
rect 1903 11512 2136 11540
rect 1903 11509 1915 11512
rect 1857 11503 1915 11509
rect 2130 11500 2136 11512
rect 2188 11500 2194 11552
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 13630 11540 13636 11552
rect 8444 11512 13636 11540
rect 8444 11500 8450 11512
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 13924 11540 13952 11648
rect 14458 11636 14464 11648
rect 14516 11676 14522 11688
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 14516 11648 15393 11676
rect 14516 11636 14522 11648
rect 15381 11645 15393 11648
rect 15427 11676 15439 11679
rect 16669 11679 16727 11685
rect 16669 11676 16681 11679
rect 15427 11648 16681 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 16669 11645 16681 11648
rect 16715 11645 16727 11679
rect 16669 11639 16727 11645
rect 14918 11540 14924 11552
rect 13924 11512 14924 11540
rect 14918 11500 14924 11512
rect 14976 11500 14982 11552
rect 15194 11540 15200 11552
rect 15155 11512 15200 11540
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 1104 11450 16468 11472
rect 1104 11398 3542 11450
rect 3594 11398 3606 11450
rect 3658 11398 3670 11450
rect 3722 11398 3734 11450
rect 3786 11398 8664 11450
rect 8716 11398 8728 11450
rect 8780 11398 8792 11450
rect 8844 11398 8856 11450
rect 8908 11398 13785 11450
rect 13837 11398 13849 11450
rect 13901 11398 13913 11450
rect 13965 11398 13977 11450
rect 14029 11398 16468 11450
rect 1104 11376 16468 11398
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 3881 11339 3939 11345
rect 3881 11336 3893 11339
rect 3476 11308 3893 11336
rect 3476 11296 3482 11308
rect 3881 11305 3893 11308
rect 3927 11305 3939 11339
rect 8386 11336 8392 11348
rect 3881 11299 3939 11305
rect 6932 11308 8392 11336
rect 3436 11268 3464 11296
rect 2976 11240 3464 11268
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11200 1731 11203
rect 1762 11200 1768 11212
rect 1719 11172 1768 11200
rect 1719 11169 1731 11172
rect 1673 11163 1731 11169
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 2130 11200 2136 11212
rect 2091 11172 2136 11200
rect 2130 11160 2136 11172
rect 2188 11160 2194 11212
rect 1486 11092 1492 11144
rect 1544 11132 1550 11144
rect 1857 11135 1915 11141
rect 1857 11132 1869 11135
rect 1544 11104 1869 11132
rect 1544 11092 1550 11104
rect 1857 11101 1869 11104
rect 1903 11101 1915 11135
rect 1857 11095 1915 11101
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11101 2007 11135
rect 1949 11095 2007 11101
rect 1964 11064 1992 11095
rect 2038 11092 2044 11144
rect 2096 11132 2102 11144
rect 2866 11132 2872 11144
rect 2096 11104 2141 11132
rect 2827 11104 2872 11132
rect 2096 11092 2102 11104
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 2976 11141 3004 11240
rect 5534 11228 5540 11280
rect 5592 11268 5598 11280
rect 6932 11268 6960 11308
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 9490 11296 9496 11348
rect 9548 11336 9554 11348
rect 11517 11339 11575 11345
rect 11517 11336 11529 11339
rect 9548 11308 11529 11336
rect 9548 11296 9554 11308
rect 11517 11305 11529 11308
rect 11563 11305 11575 11339
rect 11974 11336 11980 11348
rect 11517 11299 11575 11305
rect 11808 11308 11980 11336
rect 8018 11268 8024 11280
rect 5592 11240 6960 11268
rect 7024 11240 8024 11268
rect 5592 11228 5598 11240
rect 3145 11203 3203 11209
rect 3145 11169 3157 11203
rect 3191 11200 3203 11203
rect 3878 11200 3884 11212
rect 3191 11172 3884 11200
rect 3191 11169 3203 11172
rect 3145 11163 3203 11169
rect 3878 11160 3884 11172
rect 3936 11200 3942 11212
rect 6914 11200 6920 11212
rect 3936 11172 4200 11200
rect 3936 11160 3942 11172
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 4062 11132 4068 11144
rect 3283 11104 4068 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 4172 11141 4200 11172
rect 6288 11172 6920 11200
rect 6288 11141 6316 11172
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4433 11135 4491 11141
rect 4433 11132 4445 11135
rect 4203 11104 4445 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4433 11101 4445 11104
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 6273 11135 6331 11141
rect 6273 11101 6285 11135
rect 6319 11101 6331 11135
rect 6273 11095 6331 11101
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 7024 11132 7052 11240
rect 8018 11228 8024 11240
rect 8076 11228 8082 11280
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 7432 11172 7573 11200
rect 7432 11160 7438 11172
rect 7561 11169 7573 11172
rect 7607 11200 7619 11203
rect 8389 11203 8447 11209
rect 8389 11200 8401 11203
rect 7607 11172 8401 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 8389 11169 8401 11172
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11200 9735 11203
rect 10686 11200 10692 11212
rect 9723 11172 10692 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 6503 11104 7052 11132
rect 7285 11135 7343 11141
rect 7102 11113 7160 11119
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 2685 11067 2743 11073
rect 1964 11036 2636 11064
rect 2608 10996 2636 11036
rect 2685 11033 2697 11067
rect 2731 11064 2743 11067
rect 4080 11064 4108 11092
rect 7102 11079 7114 11113
rect 7148 11079 7160 11113
rect 7285 11101 7297 11135
rect 7331 11132 7343 11135
rect 8213 11135 8271 11141
rect 7331 11104 8156 11132
rect 7331 11101 7343 11104
rect 7285 11095 7343 11101
rect 7102 11076 7160 11079
rect 7576 11076 7604 11104
rect 4525 11067 4583 11073
rect 4525 11064 4537 11067
rect 2731 11036 2912 11064
rect 4080 11036 4537 11064
rect 2731 11033 2743 11036
rect 2685 11027 2743 11033
rect 2884 11008 2912 11036
rect 4525 11033 4537 11036
rect 4571 11033 4583 11067
rect 4525 11027 4583 11033
rect 4614 11024 4620 11076
rect 4672 11064 4678 11076
rect 6365 11067 6423 11073
rect 4672 11036 6316 11064
rect 4672 11024 4678 11036
rect 2774 10996 2780 11008
rect 2608 10968 2780 10996
rect 2774 10956 2780 10968
rect 2832 10956 2838 11008
rect 2866 10956 2872 11008
rect 2924 10956 2930 11008
rect 6288 10996 6316 11036
rect 6365 11033 6377 11067
rect 6411 11064 6423 11067
rect 6822 11064 6828 11076
rect 6411 11036 6828 11064
rect 6411 11033 6423 11036
rect 6365 11027 6423 11033
rect 6822 11024 6828 11036
rect 6880 11024 6886 11076
rect 7098 11024 7104 11076
rect 7156 11024 7162 11076
rect 7193 11067 7251 11073
rect 7193 11033 7205 11067
rect 7239 11064 7251 11067
rect 7239 11036 7328 11064
rect 7239 11033 7251 11036
rect 7193 11027 7251 11033
rect 6917 10999 6975 11005
rect 6917 10996 6929 10999
rect 6288 10968 6929 10996
rect 6917 10965 6929 10968
rect 6963 10965 6975 10999
rect 7300 10996 7328 11036
rect 7374 11024 7380 11076
rect 7432 11073 7438 11076
rect 7432 11067 7461 11073
rect 7449 11033 7461 11067
rect 7432 11027 7461 11033
rect 7432 11024 7438 11027
rect 7558 11024 7564 11076
rect 7616 11024 7622 11076
rect 8021 11067 8079 11073
rect 8021 11033 8033 11067
rect 8067 11033 8079 11067
rect 8128 11064 8156 11104
rect 8213 11101 8225 11135
rect 8259 11132 8271 11135
rect 8478 11132 8484 11144
rect 8259 11104 8484 11132
rect 8259 11101 8271 11104
rect 8213 11095 8271 11101
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 9490 11092 9496 11144
rect 9548 11132 9554 11144
rect 9585 11135 9643 11141
rect 9585 11132 9597 11135
rect 9548 11104 9597 11132
rect 9548 11092 9554 11104
rect 9585 11101 9597 11104
rect 9631 11101 9643 11135
rect 9585 11095 9643 11101
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 8128 11036 9628 11064
rect 8021 11027 8079 11033
rect 7650 10996 7656 11008
rect 7300 10968 7656 10996
rect 6917 10959 6975 10965
rect 7650 10956 7656 10968
rect 7708 10956 7714 11008
rect 8036 10996 8064 11027
rect 8202 10996 8208 11008
rect 8036 10968 8208 10996
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 8386 10956 8392 11008
rect 8444 10996 8450 11008
rect 9401 10999 9459 11005
rect 9401 10996 9413 10999
rect 8444 10968 9413 10996
rect 8444 10956 8450 10968
rect 9401 10965 9413 10968
rect 9447 10965 9459 10999
rect 9600 10996 9628 11036
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 9784 11064 9812 11095
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 10594 11132 10600 11144
rect 9916 11104 9961 11132
rect 10555 11104 10600 11132
rect 9916 11092 9922 11104
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 11808 11141 11836 11308
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 12986 11336 12992 11348
rect 12124 11308 12992 11336
rect 12124 11296 12130 11308
rect 12986 11296 12992 11308
rect 13044 11336 13050 11348
rect 13538 11336 13544 11348
rect 13044 11308 13544 11336
rect 13044 11296 13050 11308
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 13630 11296 13636 11348
rect 13688 11336 13694 11348
rect 15381 11339 15439 11345
rect 15381 11336 15393 11339
rect 13688 11308 15393 11336
rect 13688 11296 13694 11308
rect 15381 11305 15393 11308
rect 15427 11305 15439 11339
rect 15381 11299 15439 11305
rect 11882 11228 11888 11280
rect 11940 11268 11946 11280
rect 13357 11271 13415 11277
rect 13357 11268 13369 11271
rect 11940 11240 13369 11268
rect 11940 11228 11946 11240
rect 13357 11237 13369 11240
rect 13403 11237 13415 11271
rect 13357 11231 13415 11237
rect 11977 11203 12035 11209
rect 11977 11169 11989 11203
rect 12023 11200 12035 11203
rect 12621 11203 12679 11209
rect 12621 11200 12633 11203
rect 12023 11172 12633 11200
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 12621 11169 12633 11172
rect 12667 11200 12679 11203
rect 12667 11172 13216 11200
rect 12667 11169 12679 11172
rect 12621 11163 12679 11169
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11101 11759 11135
rect 11701 11095 11759 11101
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11101 12127 11135
rect 12069 11095 12127 11101
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11132 12771 11135
rect 12802 11132 12808 11144
rect 12759 11104 12808 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 9732 11036 9812 11064
rect 11716 11064 11744 11095
rect 12084 11064 12112 11095
rect 12802 11092 12808 11104
rect 12860 11092 12866 11144
rect 13188 11141 13216 11172
rect 13173 11135 13231 11141
rect 13173 11101 13185 11135
rect 13219 11101 13231 11135
rect 13372 11132 13400 11231
rect 14182 11160 14188 11212
rect 14240 11200 14246 11212
rect 14369 11203 14427 11209
rect 14369 11200 14381 11203
rect 14240 11172 14381 11200
rect 14240 11160 14246 11172
rect 14369 11169 14381 11172
rect 14415 11169 14427 11203
rect 14369 11163 14427 11169
rect 14090 11132 14096 11144
rect 13372 11104 14096 11132
rect 13173 11095 13231 11101
rect 14090 11092 14096 11104
rect 14148 11092 14154 11144
rect 15470 11092 15476 11144
rect 15528 11132 15534 11144
rect 15565 11135 15623 11141
rect 15565 11132 15577 11135
rect 15528 11104 15577 11132
rect 15528 11092 15534 11104
rect 15565 11101 15577 11104
rect 15611 11101 15623 11135
rect 15746 11132 15752 11144
rect 15707 11104 15752 11132
rect 15565 11095 15623 11101
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 12434 11064 12440 11076
rect 11716 11036 12020 11064
rect 12084 11036 12440 11064
rect 9732 11024 9738 11036
rect 10042 10996 10048 11008
rect 9600 10968 10048 10996
rect 9401 10959 9459 10965
rect 10042 10956 10048 10968
rect 10100 10956 10106 11008
rect 10318 10956 10324 11008
rect 10376 10996 10382 11008
rect 10413 10999 10471 11005
rect 10413 10996 10425 10999
rect 10376 10968 10425 10996
rect 10376 10956 10382 10968
rect 10413 10965 10425 10968
rect 10459 10965 10471 10999
rect 11992 10996 12020 11036
rect 12434 11024 12440 11036
rect 12492 11064 12498 11076
rect 12618 11064 12624 11076
rect 12492 11036 12624 11064
rect 12492 11024 12498 11036
rect 12618 11024 12624 11036
rect 12676 11024 12682 11076
rect 13354 11064 13360 11076
rect 12728 11036 13360 11064
rect 12526 10996 12532 11008
rect 11992 10968 12532 10996
rect 10413 10959 10471 10965
rect 12526 10956 12532 10968
rect 12584 10996 12590 11008
rect 12728 10996 12756 11036
rect 13354 11024 13360 11036
rect 13412 11024 13418 11076
rect 12584 10968 12756 10996
rect 12584 10956 12590 10968
rect 1104 10906 16468 10928
rect 1104 10854 6103 10906
rect 6155 10854 6167 10906
rect 6219 10854 6231 10906
rect 6283 10854 6295 10906
rect 6347 10854 11224 10906
rect 11276 10854 11288 10906
rect 11340 10854 11352 10906
rect 11404 10854 11416 10906
rect 11468 10854 16468 10906
rect 1104 10832 16468 10854
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 3878 10792 3884 10804
rect 2832 10764 2877 10792
rect 3839 10764 3884 10792
rect 2832 10752 2838 10764
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 4614 10792 4620 10804
rect 4080 10764 4620 10792
rect 1946 10684 1952 10736
rect 2004 10724 2010 10736
rect 2004 10696 2176 10724
rect 2004 10684 2010 10696
rect 2148 10665 2176 10696
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10625 2191 10659
rect 2133 10619 2191 10625
rect 2222 10616 2228 10668
rect 2280 10656 2286 10668
rect 2280 10628 2325 10656
rect 2280 10616 2286 10628
rect 2406 10616 2412 10668
rect 2464 10656 2470 10668
rect 4080 10665 4108 10764
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 4893 10795 4951 10801
rect 4893 10761 4905 10795
rect 4939 10761 4951 10795
rect 4893 10755 4951 10761
rect 6549 10795 6607 10801
rect 6549 10761 6561 10795
rect 6595 10792 6607 10795
rect 7374 10792 7380 10804
rect 6595 10764 7380 10792
rect 6595 10761 6607 10764
rect 6549 10755 6607 10761
rect 4522 10724 4528 10736
rect 4172 10696 4528 10724
rect 4172 10665 4200 10696
rect 4522 10684 4528 10696
rect 4580 10724 4586 10736
rect 4908 10724 4936 10755
rect 7374 10752 7380 10764
rect 7432 10752 7438 10804
rect 7466 10752 7472 10804
rect 7524 10792 7530 10804
rect 8202 10792 8208 10804
rect 7524 10764 8208 10792
rect 7524 10752 7530 10764
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 10689 10795 10747 10801
rect 10689 10792 10701 10795
rect 10468 10764 10701 10792
rect 10468 10752 10474 10764
rect 10689 10761 10701 10764
rect 10735 10761 10747 10795
rect 10962 10792 10968 10804
rect 10923 10764 10968 10792
rect 10689 10755 10747 10761
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 11882 10792 11888 10804
rect 11716 10764 11888 10792
rect 4580 10696 4936 10724
rect 4580 10684 4586 10696
rect 9398 10684 9404 10736
rect 9456 10724 9462 10736
rect 11716 10733 11744 10764
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 13265 10795 13323 10801
rect 13265 10761 13277 10795
rect 13311 10792 13323 10795
rect 14274 10792 14280 10804
rect 13311 10764 14280 10792
rect 13311 10761 13323 10764
rect 13265 10755 13323 10761
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 15470 10792 15476 10804
rect 15431 10764 15476 10792
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 9585 10727 9643 10733
rect 9585 10724 9597 10727
rect 9456 10696 9597 10724
rect 9456 10684 9462 10696
rect 9585 10693 9597 10696
rect 9631 10693 9643 10727
rect 9585 10687 9643 10693
rect 9815 10727 9873 10733
rect 9815 10693 9827 10727
rect 9861 10724 9873 10727
rect 11517 10727 11575 10733
rect 11517 10724 11529 10727
rect 9861 10696 11529 10724
rect 9861 10693 9873 10696
rect 9815 10687 9873 10693
rect 11517 10693 11529 10696
rect 11563 10693 11575 10727
rect 11517 10687 11575 10693
rect 11701 10727 11759 10733
rect 11701 10693 11713 10727
rect 11747 10693 11759 10727
rect 11701 10687 11759 10693
rect 11790 10684 11796 10736
rect 11848 10724 11854 10736
rect 12897 10727 12955 10733
rect 12897 10724 12909 10727
rect 11848 10696 12909 10724
rect 11848 10684 11854 10696
rect 12897 10693 12909 10696
rect 12943 10693 12955 10727
rect 12897 10687 12955 10693
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 2464 10628 2697 10656
rect 2464 10616 2470 10628
rect 2685 10625 2697 10628
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10656 4491 10659
rect 4890 10656 4896 10668
rect 4479 10628 4896 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5169 10659 5227 10665
rect 5169 10656 5181 10659
rect 5000 10628 5181 10656
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10588 2007 10591
rect 3234 10588 3240 10600
rect 1995 10560 3240 10588
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10588 4399 10591
rect 5000 10588 5028 10628
rect 5169 10625 5181 10628
rect 5215 10656 5227 10659
rect 5442 10656 5448 10668
rect 5215 10628 5448 10656
rect 5215 10625 5227 10628
rect 5169 10619 5227 10625
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 7098 10656 7104 10668
rect 6687 10628 7104 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10656 7343 10659
rect 8386 10656 8392 10668
rect 7331 10628 8392 10656
rect 7331 10625 7343 10628
rect 7285 10619 7343 10625
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 9490 10656 9496 10668
rect 9451 10628 9496 10656
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 9732 10628 9825 10656
rect 9732 10616 9738 10628
rect 10042 10616 10048 10668
rect 10100 10656 10106 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 10100 10628 10609 10656
rect 10100 10616 10106 10628
rect 10597 10625 10609 10628
rect 10643 10625 10655 10659
rect 10597 10619 10655 10625
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10656 10839 10659
rect 10827 10628 11008 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 4387 10560 5028 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 5132 10560 5549 10588
rect 5132 10548 5138 10560
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 5537 10551 5595 10557
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 7742 10588 7748 10600
rect 7432 10560 7748 10588
rect 7432 10548 7438 10560
rect 7742 10548 7748 10560
rect 7800 10548 7806 10600
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10588 8079 10591
rect 8110 10588 8116 10600
rect 8067 10560 8116 10588
rect 8067 10557 8079 10560
rect 8021 10551 8079 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 9122 10548 9128 10600
rect 9180 10588 9186 10600
rect 9692 10588 9720 10616
rect 9950 10588 9956 10600
rect 9180 10560 9720 10588
rect 9911 10560 9956 10588
rect 9180 10548 9186 10560
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 10612 10588 10640 10619
rect 10870 10588 10876 10600
rect 10244 10560 10548 10588
rect 10612 10560 10876 10588
rect 5626 10480 5632 10532
rect 5684 10520 5690 10532
rect 9309 10523 9367 10529
rect 9309 10520 9321 10523
rect 5684 10492 9321 10520
rect 5684 10480 5690 10492
rect 9309 10489 9321 10492
rect 9355 10489 9367 10523
rect 10244 10520 10272 10560
rect 9309 10483 9367 10489
rect 9646 10492 10272 10520
rect 1854 10412 1860 10464
rect 1912 10452 1918 10464
rect 2041 10455 2099 10461
rect 2041 10452 2053 10455
rect 1912 10424 2053 10452
rect 1912 10412 1918 10424
rect 2041 10421 2053 10424
rect 2087 10421 2099 10455
rect 7190 10452 7196 10464
rect 7103 10424 7196 10452
rect 2041 10415 2099 10421
rect 7190 10412 7196 10424
rect 7248 10452 7254 10464
rect 7742 10452 7748 10464
rect 7248 10424 7748 10452
rect 7248 10412 7254 10424
rect 7742 10412 7748 10424
rect 7800 10412 7806 10464
rect 9030 10412 9036 10464
rect 9088 10452 9094 10464
rect 9646 10452 9674 10492
rect 10318 10480 10324 10532
rect 10376 10520 10382 10532
rect 10413 10523 10471 10529
rect 10413 10520 10425 10523
rect 10376 10492 10425 10520
rect 10376 10480 10382 10492
rect 10413 10489 10425 10492
rect 10459 10489 10471 10523
rect 10520 10520 10548 10560
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 10980 10588 11008 10628
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11882 10656 11888 10668
rect 11112 10628 11888 10656
rect 11112 10616 11118 10628
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 12713 10659 12771 10665
rect 12713 10656 12725 10659
rect 12492 10628 12725 10656
rect 12492 10616 12498 10628
rect 12713 10625 12725 10628
rect 12759 10625 12771 10659
rect 12986 10656 12992 10668
rect 12947 10628 12992 10656
rect 12713 10619 12771 10625
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 13909 10659 13967 10665
rect 13909 10625 13921 10659
rect 13955 10656 13967 10659
rect 14366 10656 14372 10668
rect 13955 10628 14372 10656
rect 13955 10625 13967 10628
rect 13909 10619 13967 10625
rect 12802 10588 12808 10600
rect 10980 10560 12808 10588
rect 10980 10520 11008 10560
rect 12802 10548 12808 10560
rect 12860 10588 12866 10600
rect 13096 10588 13124 10619
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 14918 10656 14924 10668
rect 14879 10628 14924 10656
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 15102 10616 15108 10668
rect 15160 10656 15166 10668
rect 15197 10659 15255 10665
rect 15197 10656 15209 10659
rect 15160 10628 15209 10656
rect 15160 10616 15166 10628
rect 15197 10625 15209 10628
rect 15243 10625 15255 10659
rect 15197 10619 15255 10625
rect 15289 10659 15347 10665
rect 15289 10625 15301 10659
rect 15335 10656 15347 10659
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 15335 10628 16681 10656
rect 15335 10625 15347 10628
rect 15289 10619 15347 10625
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 12860 10560 13124 10588
rect 12860 10548 12866 10560
rect 10520 10492 11008 10520
rect 10413 10483 10471 10489
rect 13538 10480 13544 10532
rect 13596 10520 13602 10532
rect 13725 10523 13783 10529
rect 13725 10520 13737 10523
rect 13596 10492 13737 10520
rect 13596 10480 13602 10492
rect 13725 10489 13737 10492
rect 13771 10520 13783 10523
rect 15013 10523 15071 10529
rect 15013 10520 15025 10523
rect 13771 10492 15025 10520
rect 13771 10489 13783 10492
rect 13725 10483 13783 10489
rect 15013 10489 15025 10492
rect 15059 10520 15071 10523
rect 15194 10520 15200 10532
rect 15059 10492 15200 10520
rect 15059 10489 15071 10492
rect 15013 10483 15071 10489
rect 15194 10480 15200 10492
rect 15252 10480 15258 10532
rect 9088 10424 9674 10452
rect 9088 10412 9094 10424
rect 10134 10412 10140 10464
rect 10192 10452 10198 10464
rect 11790 10452 11796 10464
rect 10192 10424 11796 10452
rect 10192 10412 10198 10424
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 1104 10362 16468 10384
rect 1104 10310 3542 10362
rect 3594 10310 3606 10362
rect 3658 10310 3670 10362
rect 3722 10310 3734 10362
rect 3786 10310 8664 10362
rect 8716 10310 8728 10362
rect 8780 10310 8792 10362
rect 8844 10310 8856 10362
rect 8908 10310 13785 10362
rect 13837 10310 13849 10362
rect 13901 10310 13913 10362
rect 13965 10310 13977 10362
rect 14029 10310 16468 10362
rect 1104 10288 16468 10310
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 2593 10251 2651 10257
rect 2593 10248 2605 10251
rect 2280 10220 2605 10248
rect 2280 10208 2286 10220
rect 2593 10217 2605 10220
rect 2639 10217 2651 10251
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 2593 10211 2651 10217
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 7098 10208 7104 10260
rect 7156 10248 7162 10260
rect 7745 10251 7803 10257
rect 7745 10248 7757 10251
rect 7156 10220 7757 10248
rect 7156 10208 7162 10220
rect 7745 10217 7757 10220
rect 7791 10217 7803 10251
rect 9766 10248 9772 10260
rect 9727 10220 9772 10248
rect 7745 10211 7803 10217
rect 9766 10208 9772 10220
rect 9824 10208 9830 10260
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 10778 10248 10784 10260
rect 10008 10220 10784 10248
rect 10008 10208 10014 10220
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 10870 10208 10876 10260
rect 10928 10248 10934 10260
rect 10928 10220 11468 10248
rect 10928 10208 10934 10220
rect 2866 10180 2872 10192
rect 2792 10152 2872 10180
rect 1489 10115 1547 10121
rect 1489 10081 1501 10115
rect 1535 10112 1547 10115
rect 1946 10112 1952 10124
rect 1535 10084 1952 10112
rect 1535 10081 1547 10084
rect 1489 10075 1547 10081
rect 1946 10072 1952 10084
rect 2004 10112 2010 10124
rect 2406 10112 2412 10124
rect 2004 10084 2412 10112
rect 2004 10072 2010 10084
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 2792 10121 2820 10152
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 6822 10140 6828 10192
rect 6880 10180 6886 10192
rect 6880 10152 8248 10180
rect 6880 10140 6886 10152
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10112 2835 10115
rect 5902 10112 5908 10124
rect 2823 10084 3832 10112
rect 5863 10084 5908 10112
rect 2823 10081 2835 10084
rect 2777 10075 2835 10081
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 1854 10044 1860 10056
rect 1627 10016 1860 10044
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 1854 10004 1860 10016
rect 1912 10004 1918 10056
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10044 2927 10047
rect 3050 10044 3056 10056
rect 2915 10016 3056 10044
rect 2915 10013 2927 10016
rect 2869 10007 2927 10013
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 3234 10044 3240 10056
rect 3195 10016 3240 10044
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 3804 10053 3832 10084
rect 5902 10072 5908 10084
rect 5960 10072 5966 10124
rect 8018 10112 8024 10124
rect 7979 10084 8024 10112
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8220 10121 8248 10152
rect 9674 10140 9680 10192
rect 9732 10180 9738 10192
rect 11440 10180 11468 10220
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 12069 10251 12127 10257
rect 12069 10248 12081 10251
rect 12032 10220 12081 10248
rect 12032 10208 12038 10220
rect 12069 10217 12081 10220
rect 12115 10217 12127 10251
rect 12069 10211 12127 10217
rect 13265 10251 13323 10257
rect 13265 10217 13277 10251
rect 13311 10248 13323 10251
rect 16577 10251 16635 10257
rect 16577 10248 16589 10251
rect 13311 10220 16589 10248
rect 13311 10217 13323 10220
rect 13265 10211 13323 10217
rect 16577 10217 16589 10220
rect 16623 10217 16635 10251
rect 16577 10211 16635 10217
rect 13078 10180 13084 10192
rect 9732 10152 11284 10180
rect 11440 10152 13084 10180
rect 9732 10140 9738 10152
rect 8205 10115 8263 10121
rect 8205 10081 8217 10115
rect 8251 10081 8263 10115
rect 8205 10075 8263 10081
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 5626 10044 5632 10056
rect 5587 10016 5632 10044
rect 3789 10007 3847 10013
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 5718 10004 5724 10056
rect 5776 10044 5782 10056
rect 5997 10047 6055 10053
rect 5776 10016 5821 10044
rect 5776 10004 5782 10016
rect 5997 10013 6009 10047
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10044 7159 10047
rect 7926 10044 7932 10056
rect 7147 10016 7932 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 3068 9976 3096 10004
rect 3973 9979 4031 9985
rect 3973 9976 3985 9979
rect 3068 9948 3985 9976
rect 3973 9945 3985 9948
rect 4019 9945 4031 9979
rect 3973 9939 4031 9945
rect 5810 9936 5816 9988
rect 5868 9976 5874 9988
rect 6012 9976 6040 10007
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 8122 10047 8180 10053
rect 8122 10013 8134 10047
rect 8168 10044 8180 10047
rect 8386 10044 8392 10056
rect 8168 10016 8248 10044
rect 8347 10016 8392 10044
rect 8168 10013 8180 10016
rect 8122 10007 8180 10013
rect 5868 9948 6040 9976
rect 6917 9979 6975 9985
rect 5868 9936 5874 9948
rect 6917 9945 6929 9979
rect 6963 9976 6975 9979
rect 7466 9976 7472 9988
rect 6963 9948 7472 9976
rect 6963 9945 6975 9948
rect 6917 9939 6975 9945
rect 7466 9936 7472 9948
rect 7524 9936 7530 9988
rect 7742 9936 7748 9988
rect 7800 9976 7806 9988
rect 8220 9976 8248 10016
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10044 8999 10047
rect 9030 10044 9036 10056
rect 8987 10016 9036 10044
rect 8987 10013 8999 10016
rect 8941 10007 8999 10013
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 10152 10053 10180 10152
rect 10318 10112 10324 10124
rect 10279 10084 10324 10112
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 10778 10072 10784 10124
rect 10836 10112 10842 10124
rect 11149 10115 11207 10121
rect 11149 10112 11161 10115
rect 10836 10084 11161 10112
rect 10836 10072 10842 10084
rect 11149 10081 11161 10084
rect 11195 10081 11207 10115
rect 11149 10075 11207 10081
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 7800 9948 8248 9976
rect 7800 9936 7806 9948
rect 9858 9936 9864 9988
rect 9916 9976 9922 9988
rect 10781 9979 10839 9985
rect 9916 9948 10364 9976
rect 9916 9936 9922 9948
rect 2038 9868 2044 9920
rect 2096 9908 2102 9920
rect 2133 9911 2191 9917
rect 2133 9908 2145 9911
rect 2096 9880 2145 9908
rect 2096 9868 2102 9880
rect 2133 9877 2145 9880
rect 2179 9877 2191 9911
rect 2133 9871 2191 9877
rect 3234 9868 3240 9920
rect 3292 9908 3298 9920
rect 4157 9911 4215 9917
rect 4157 9908 4169 9911
rect 3292 9880 4169 9908
rect 3292 9868 3298 9880
rect 4157 9877 4169 9880
rect 4203 9877 4215 9911
rect 4157 9871 4215 9877
rect 7285 9911 7343 9917
rect 7285 9877 7297 9911
rect 7331 9908 7343 9911
rect 7558 9908 7564 9920
rect 7331 9880 7564 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 7558 9868 7564 9880
rect 7616 9868 7622 9920
rect 9122 9908 9128 9920
rect 9083 9880 9128 9908
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 9953 9911 10011 9917
rect 9953 9908 9965 9911
rect 9732 9880 9965 9908
rect 9732 9868 9738 9880
rect 9953 9877 9965 9880
rect 9999 9877 10011 9911
rect 9953 9871 10011 9877
rect 10045 9911 10103 9917
rect 10045 9877 10057 9911
rect 10091 9908 10103 9911
rect 10134 9908 10140 9920
rect 10091 9880 10140 9908
rect 10091 9877 10103 9880
rect 10045 9871 10103 9877
rect 10134 9868 10140 9880
rect 10192 9868 10198 9920
rect 10336 9908 10364 9948
rect 10781 9945 10793 9979
rect 10827 9945 10839 9979
rect 10781 9939 10839 9945
rect 10965 9979 11023 9985
rect 10965 9945 10977 9979
rect 11011 9976 11023 9979
rect 11054 9976 11060 9988
rect 11011 9948 11060 9976
rect 11011 9945 11023 9948
rect 10965 9939 11023 9945
rect 10796 9908 10824 9939
rect 11054 9936 11060 9948
rect 11112 9936 11118 9988
rect 10336 9880 10824 9908
rect 11256 9908 11284 10152
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 14918 10072 14924 10124
rect 14976 10112 14982 10124
rect 15381 10115 15439 10121
rect 15381 10112 15393 10115
rect 14976 10084 15393 10112
rect 14976 10072 14982 10084
rect 15381 10081 15393 10084
rect 15427 10081 15439 10115
rect 15381 10075 15439 10081
rect 13078 10044 13084 10056
rect 13039 10016 13084 10044
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 14090 10044 14096 10056
rect 14051 10016 14096 10044
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 15102 10044 15108 10056
rect 15063 10016 15108 10044
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 11974 9976 11980 9988
rect 11935 9948 11980 9976
rect 11974 9936 11980 9948
rect 12032 9936 12038 9988
rect 12434 9936 12440 9988
rect 12492 9976 12498 9988
rect 12618 9976 12624 9988
rect 12492 9948 12624 9976
rect 12492 9936 12498 9948
rect 12618 9936 12624 9948
rect 12676 9976 12682 9988
rect 12713 9979 12771 9985
rect 12713 9976 12725 9979
rect 12676 9948 12725 9976
rect 12676 9936 12682 9948
rect 12713 9945 12725 9948
rect 12759 9945 12771 9979
rect 12713 9939 12771 9945
rect 14182 9936 14188 9988
rect 14240 9976 14246 9988
rect 14277 9979 14335 9985
rect 14277 9976 14289 9979
rect 14240 9948 14289 9976
rect 14240 9936 14246 9948
rect 14277 9945 14289 9948
rect 14323 9976 14335 9979
rect 14642 9976 14648 9988
rect 14323 9948 14648 9976
rect 14323 9945 14335 9948
rect 14277 9939 14335 9945
rect 14642 9936 14648 9948
rect 14700 9936 14706 9988
rect 12897 9911 12955 9917
rect 12897 9908 12909 9911
rect 11256 9880 12909 9908
rect 12897 9877 12909 9880
rect 12943 9877 12955 9911
rect 12897 9871 12955 9877
rect 12986 9868 12992 9920
rect 13044 9908 13050 9920
rect 14458 9908 14464 9920
rect 13044 9880 13089 9908
rect 14419 9880 14464 9908
rect 13044 9868 13050 9880
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 1104 9818 16468 9840
rect 1104 9766 6103 9818
rect 6155 9766 6167 9818
rect 6219 9766 6231 9818
rect 6283 9766 6295 9818
rect 6347 9766 11224 9818
rect 11276 9766 11288 9818
rect 11340 9766 11352 9818
rect 11404 9766 11416 9818
rect 11468 9766 16468 9818
rect 1104 9744 16468 9766
rect 1857 9707 1915 9713
rect 1857 9673 1869 9707
rect 1903 9704 1915 9707
rect 1946 9704 1952 9716
rect 1903 9676 1952 9704
rect 1903 9673 1915 9676
rect 1857 9667 1915 9673
rect 1946 9664 1952 9676
rect 2004 9664 2010 9716
rect 7006 9664 7012 9716
rect 7064 9704 7070 9716
rect 8110 9704 8116 9716
rect 7064 9676 8116 9704
rect 7064 9664 7070 9676
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8481 9707 8539 9713
rect 8481 9673 8493 9707
rect 8527 9704 8539 9707
rect 9490 9704 9496 9716
rect 8527 9676 9496 9704
rect 8527 9673 8539 9676
rect 8481 9667 8539 9673
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 9677 9707 9735 9713
rect 9677 9673 9689 9707
rect 9723 9704 9735 9707
rect 9766 9704 9772 9716
rect 9723 9676 9772 9704
rect 9723 9673 9735 9676
rect 9677 9667 9735 9673
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 9950 9704 9956 9716
rect 9876 9676 9956 9704
rect 5721 9639 5779 9645
rect 5721 9605 5733 9639
rect 5767 9636 5779 9639
rect 5902 9636 5908 9648
rect 5767 9608 5908 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2222 9528 2228 9580
rect 2280 9568 2286 9580
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 2280 9540 2881 9568
rect 2280 9528 2286 9540
rect 2869 9537 2881 9540
rect 2915 9537 2927 9571
rect 2869 9531 2927 9537
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9568 3019 9571
rect 3234 9568 3240 9580
rect 3007 9540 3240 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 5736 9568 5764 9599
rect 5902 9596 5908 9608
rect 5960 9636 5966 9648
rect 9876 9636 9904 9676
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 5960 9608 8524 9636
rect 5960 9596 5966 9608
rect 7282 9568 7288 9580
rect 5491 9540 5764 9568
rect 7243 9540 7288 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 7558 9568 7564 9580
rect 7519 9540 7564 9568
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 7742 9568 7748 9580
rect 7703 9540 7748 9568
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 2148 9500 2176 9528
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2148 9472 2697 9500
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9500 5411 9503
rect 5810 9500 5816 9512
rect 5399 9472 5816 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 5810 9460 5816 9472
rect 5868 9460 5874 9512
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9500 7527 9503
rect 8386 9500 8392 9512
rect 7515 9472 8392 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 8496 9500 8524 9608
rect 8588 9608 9904 9636
rect 8588 9577 8616 9608
rect 8573 9571 8631 9577
rect 8573 9537 8585 9571
rect 8619 9537 8631 9571
rect 8573 9531 8631 9537
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9582 9568 9588 9580
rect 9079 9540 9588 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 9582 9528 9588 9540
rect 9640 9568 9646 9580
rect 9861 9571 9919 9577
rect 9861 9568 9873 9571
rect 9640 9540 9873 9568
rect 9640 9528 9646 9540
rect 9861 9537 9873 9540
rect 9907 9537 9919 9571
rect 9950 9552 9956 9604
rect 10008 9552 10014 9604
rect 11698 9596 11704 9648
rect 11756 9636 11762 9648
rect 12161 9639 12219 9645
rect 12161 9636 12173 9639
rect 11756 9608 12173 9636
rect 11756 9596 11762 9608
rect 12161 9605 12173 9608
rect 12207 9605 12219 9639
rect 12161 9599 12219 9605
rect 14645 9639 14703 9645
rect 14645 9605 14657 9639
rect 14691 9636 14703 9639
rect 14734 9636 14740 9648
rect 14691 9608 14740 9636
rect 14691 9605 14703 9608
rect 14645 9599 14703 9605
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 10045 9571 10103 9577
rect 9861 9531 9919 9537
rect 9953 9537 9965 9552
rect 9999 9537 10011 9552
rect 9953 9531 10011 9537
rect 10045 9537 10057 9571
rect 10091 9568 10103 9571
rect 10594 9568 10600 9580
rect 10091 9540 10600 9568
rect 10091 9537 10103 9540
rect 10045 9531 10103 9537
rect 10594 9528 10600 9540
rect 10652 9568 10658 9580
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 10652 9540 10793 9568
rect 10652 9528 10658 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9568 10931 9571
rect 11606 9568 11612 9580
rect 10919 9540 11612 9568
rect 10919 9537 10931 9540
rect 10873 9531 10931 9537
rect 11606 9528 11612 9540
rect 11664 9568 11670 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11664 9540 11805 9568
rect 11664 9528 11670 9540
rect 11793 9537 11805 9540
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 12526 9528 12532 9580
rect 12584 9568 12590 9580
rect 12894 9568 12900 9580
rect 12584 9540 12900 9568
rect 12584 9528 12590 9540
rect 12894 9528 12900 9540
rect 12952 9568 12958 9580
rect 13081 9571 13139 9577
rect 13081 9568 13093 9571
rect 12952 9540 13093 9568
rect 12952 9528 12958 9540
rect 13081 9537 13093 9540
rect 13127 9537 13139 9571
rect 13081 9531 13139 9537
rect 13538 9528 13544 9580
rect 13596 9568 13602 9580
rect 13817 9571 13875 9577
rect 13817 9568 13829 9571
rect 13596 9540 13829 9568
rect 13596 9528 13602 9540
rect 13817 9537 13829 9540
rect 13863 9568 13875 9571
rect 14093 9571 14151 9577
rect 14093 9568 14105 9571
rect 13863 9540 14105 9568
rect 13863 9537 13875 9540
rect 13817 9531 13875 9537
rect 14093 9537 14105 9540
rect 14139 9537 14151 9571
rect 14826 9568 14832 9580
rect 14787 9540 14832 9568
rect 14093 9531 14151 9537
rect 14826 9528 14832 9540
rect 14884 9528 14890 9580
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9568 15163 9571
rect 15194 9568 15200 9580
rect 15151 9540 15200 9568
rect 15151 9537 15163 9540
rect 15105 9531 15163 9537
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15286 9528 15292 9580
rect 15344 9568 15350 9580
rect 15344 9540 15389 9568
rect 15344 9528 15350 9540
rect 13725 9503 13783 9509
rect 8496 9472 13676 9500
rect 2777 9435 2835 9441
rect 2777 9401 2789 9435
rect 2823 9432 2835 9435
rect 2958 9432 2964 9444
rect 2823 9404 2964 9432
rect 2823 9401 2835 9404
rect 2777 9395 2835 9401
rect 2958 9392 2964 9404
rect 3016 9392 3022 9444
rect 7190 9392 7196 9444
rect 7248 9432 7254 9444
rect 7377 9435 7435 9441
rect 7377 9432 7389 9435
rect 7248 9404 7389 9432
rect 7248 9392 7254 9404
rect 7377 9401 7389 9404
rect 7423 9401 7435 9435
rect 7377 9395 7435 9401
rect 8294 9392 8300 9444
rect 8352 9432 8358 9444
rect 10229 9435 10287 9441
rect 10229 9432 10241 9435
rect 8352 9404 10241 9432
rect 8352 9392 8358 9404
rect 10229 9401 10241 9404
rect 10275 9432 10287 9435
rect 13078 9432 13084 9444
rect 10275 9404 13084 9432
rect 10275 9401 10287 9404
rect 10229 9395 10287 9401
rect 13078 9392 13084 9404
rect 13136 9392 13142 9444
rect 13446 9392 13452 9444
rect 13504 9432 13510 9444
rect 13541 9435 13599 9441
rect 13541 9432 13553 9435
rect 13504 9404 13553 9432
rect 13504 9392 13510 9404
rect 13541 9401 13553 9404
rect 13587 9401 13599 9435
rect 13541 9395 13599 9401
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5718 9364 5724 9376
rect 5215 9336 5724 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 7101 9367 7159 9373
rect 7101 9364 7113 9367
rect 6052 9336 7113 9364
rect 6052 9324 6058 9336
rect 7101 9333 7113 9336
rect 7147 9333 7159 9367
rect 7101 9327 7159 9333
rect 9217 9367 9275 9373
rect 9217 9333 9229 9367
rect 9263 9364 9275 9367
rect 9674 9364 9680 9376
rect 9263 9336 9680 9364
rect 9263 9333 9275 9336
rect 9217 9327 9275 9333
rect 9674 9324 9680 9336
rect 9732 9364 9738 9376
rect 10502 9364 10508 9376
rect 9732 9336 10508 9364
rect 9732 9324 9738 9336
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 12897 9367 12955 9373
rect 12897 9364 12909 9367
rect 12768 9336 12909 9364
rect 12768 9324 12774 9336
rect 12897 9333 12909 9336
rect 12943 9333 12955 9367
rect 13648 9364 13676 9472
rect 13725 9469 13737 9503
rect 13771 9500 13783 9503
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 13771 9472 14197 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 14185 9469 14197 9472
rect 14231 9500 14243 9503
rect 14458 9500 14464 9512
rect 14231 9472 14464 9500
rect 14231 9469 14243 9472
rect 14185 9463 14243 9469
rect 14458 9460 14464 9472
rect 14516 9500 14522 9512
rect 14734 9500 14740 9512
rect 14516 9472 14740 9500
rect 14516 9460 14522 9472
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 14458 9364 14464 9376
rect 13648 9336 14464 9364
rect 12897 9327 12955 9333
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 1104 9274 16468 9296
rect 1104 9222 3542 9274
rect 3594 9222 3606 9274
rect 3658 9222 3670 9274
rect 3722 9222 3734 9274
rect 3786 9222 8664 9274
rect 8716 9222 8728 9274
rect 8780 9222 8792 9274
rect 8844 9222 8856 9274
rect 8908 9222 13785 9274
rect 13837 9222 13849 9274
rect 13901 9222 13913 9274
rect 13965 9222 13977 9274
rect 14029 9222 16468 9274
rect 1104 9200 16468 9222
rect 2130 9160 2136 9172
rect 2091 9132 2136 9160
rect 2130 9120 2136 9132
rect 2188 9120 2194 9172
rect 3881 9163 3939 9169
rect 3881 9129 3893 9163
rect 3927 9160 3939 9163
rect 4062 9160 4068 9172
rect 3927 9132 4068 9160
rect 3927 9129 3939 9132
rect 3881 9123 3939 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 10226 9160 10232 9172
rect 5736 9132 10232 9160
rect 5736 9092 5764 9132
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 11054 9120 11060 9172
rect 11112 9160 11118 9172
rect 11149 9163 11207 9169
rect 11149 9160 11161 9163
rect 11112 9132 11161 9160
rect 11112 9120 11118 9132
rect 11149 9129 11161 9132
rect 11195 9129 11207 9163
rect 11606 9160 11612 9172
rect 11567 9132 11612 9160
rect 11149 9123 11207 9129
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 13538 9160 13544 9172
rect 13499 9132 13544 9160
rect 13538 9120 13544 9132
rect 13596 9120 13602 9172
rect 14093 9163 14151 9169
rect 14093 9129 14105 9163
rect 14139 9160 14151 9163
rect 14550 9160 14556 9172
rect 14139 9132 14556 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 2792 9064 5764 9092
rect 2792 8965 2820 9064
rect 5810 9052 5816 9104
rect 5868 9092 5874 9104
rect 13446 9092 13452 9104
rect 5868 9064 13452 9092
rect 5868 9052 5874 9064
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 9024 4123 9027
rect 4338 9024 4344 9036
rect 4111 8996 4344 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 4338 8984 4344 8996
rect 4396 9024 4402 9036
rect 4525 9027 4583 9033
rect 4525 9024 4537 9027
rect 4396 8996 4537 9024
rect 4396 8984 4402 8996
rect 4525 8993 4537 8996
rect 4571 9024 4583 9027
rect 7285 9027 7343 9033
rect 7285 9024 7297 9027
rect 4571 8996 7297 9024
rect 4571 8993 4583 8996
rect 4525 8987 4583 8993
rect 7285 8993 7297 8996
rect 7331 8993 7343 9027
rect 7285 8987 7343 8993
rect 7558 8984 7564 9036
rect 7616 9024 7622 9036
rect 7929 9027 7987 9033
rect 7929 9024 7941 9027
rect 7616 8996 7941 9024
rect 7616 8984 7622 8996
rect 7929 8993 7941 8996
rect 7975 8993 7987 9027
rect 9122 9024 9128 9036
rect 7929 8987 7987 8993
rect 8220 8996 9128 9024
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8925 2835 8959
rect 2777 8919 2835 8925
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 6825 8959 6883 8965
rect 6825 8925 6837 8959
rect 6871 8956 6883 8959
rect 7466 8956 7472 8968
rect 6871 8928 7472 8956
rect 6871 8925 6883 8928
rect 6825 8919 6883 8925
rect 1765 8891 1823 8897
rect 1765 8857 1777 8891
rect 1811 8888 1823 8891
rect 1854 8888 1860 8900
rect 1811 8860 1860 8888
rect 1811 8857 1823 8860
rect 1765 8851 1823 8857
rect 1854 8848 1860 8860
rect 1912 8848 1918 8900
rect 1946 8848 1952 8900
rect 2004 8888 2010 8900
rect 4172 8888 4200 8919
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 8220 8956 8248 8996
rect 9122 8984 9128 8996
rect 9180 8984 9186 9036
rect 9217 9027 9275 9033
rect 9217 8993 9229 9027
rect 9263 9024 9275 9027
rect 10134 9024 10140 9036
rect 9263 8996 10140 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 9024 10655 9027
rect 11974 9024 11980 9036
rect 10643 8996 11980 9024
rect 10643 8993 10655 8996
rect 10597 8987 10655 8993
rect 7699 8928 8248 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8352 8928 8953 8956
rect 8352 8916 8358 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9582 8916 9588 8968
rect 9640 8956 9646 8968
rect 11440 8965 11468 8996
rect 11974 8984 11980 8996
rect 12032 8984 12038 9036
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 13556 9024 13584 9120
rect 12492 8996 12537 9024
rect 13556 8996 14596 9024
rect 12492 8984 12498 8996
rect 10505 8959 10563 8965
rect 10505 8956 10517 8959
rect 9640 8928 10517 8956
rect 9640 8916 9646 8928
rect 10505 8925 10517 8928
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 11333 8959 11391 8965
rect 11333 8925 11345 8959
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8925 11759 8959
rect 11701 8919 11759 8925
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8956 13415 8959
rect 14090 8956 14096 8968
rect 13403 8928 14096 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 4430 8888 4436 8900
rect 2004 8860 2049 8888
rect 4172 8860 4436 8888
rect 2004 8848 2010 8860
rect 4430 8848 4436 8860
rect 4488 8848 4494 8900
rect 6733 8891 6791 8897
rect 6733 8857 6745 8891
rect 6779 8888 6791 8891
rect 6779 8860 7512 8888
rect 6779 8857 6791 8860
rect 6733 8851 6791 8857
rect 2685 8823 2743 8829
rect 2685 8789 2697 8823
rect 2731 8820 2743 8823
rect 2866 8820 2872 8832
rect 2731 8792 2872 8820
rect 2731 8789 2743 8792
rect 2685 8783 2743 8789
rect 2866 8780 2872 8792
rect 2924 8780 2930 8832
rect 7484 8820 7512 8860
rect 7558 8848 7564 8900
rect 7616 8888 7622 8900
rect 7616 8860 7661 8888
rect 7616 8848 7622 8860
rect 7742 8848 7748 8900
rect 7800 8897 7806 8900
rect 7800 8891 7829 8897
rect 7817 8888 7829 8891
rect 11348 8888 11376 8919
rect 11514 8888 11520 8900
rect 7817 8860 7893 8888
rect 11348 8860 11520 8888
rect 7817 8857 7829 8860
rect 7800 8851 7829 8857
rect 7800 8848 7806 8851
rect 11514 8848 11520 8860
rect 11572 8848 11578 8900
rect 11716 8888 11744 8919
rect 14090 8916 14096 8928
rect 14148 8916 14154 8968
rect 14568 8965 14596 8996
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14734 8956 14740 8968
rect 14695 8928 14740 8956
rect 14553 8919 14611 8925
rect 12253 8891 12311 8897
rect 12253 8888 12265 8891
rect 11716 8860 12265 8888
rect 12253 8857 12265 8860
rect 12299 8888 12311 8891
rect 12342 8888 12348 8900
rect 12299 8860 12348 8888
rect 12299 8857 12311 8860
rect 12253 8851 12311 8857
rect 12342 8848 12348 8860
rect 12400 8848 12406 8900
rect 13173 8891 13231 8897
rect 13173 8857 13185 8891
rect 13219 8888 13231 8891
rect 13446 8888 13452 8900
rect 13219 8860 13452 8888
rect 13219 8857 13231 8860
rect 13173 8851 13231 8857
rect 13446 8848 13452 8860
rect 13504 8888 13510 8900
rect 14292 8888 14320 8919
rect 14734 8916 14740 8928
rect 14792 8916 14798 8968
rect 13504 8860 14320 8888
rect 13504 8848 13510 8860
rect 14918 8848 14924 8900
rect 14976 8888 14982 8900
rect 15473 8891 15531 8897
rect 15473 8888 15485 8891
rect 14976 8860 15485 8888
rect 14976 8848 14982 8860
rect 15473 8857 15485 8860
rect 15519 8857 15531 8891
rect 15654 8888 15660 8900
rect 15615 8860 15660 8888
rect 15473 8851 15531 8857
rect 15654 8848 15660 8860
rect 15712 8848 15718 8900
rect 7760 8820 7788 8848
rect 7484 8792 7788 8820
rect 1104 8730 16468 8752
rect 1104 8678 6103 8730
rect 6155 8678 6167 8730
rect 6219 8678 6231 8730
rect 6283 8678 6295 8730
rect 6347 8678 11224 8730
rect 11276 8678 11288 8730
rect 11340 8678 11352 8730
rect 11404 8678 11416 8730
rect 11468 8678 16468 8730
rect 1104 8656 16468 8678
rect 1673 8619 1731 8625
rect 1673 8585 1685 8619
rect 1719 8616 1731 8619
rect 2222 8616 2228 8628
rect 1719 8588 2228 8616
rect 1719 8585 1731 8588
rect 1673 8579 1731 8585
rect 2222 8576 2228 8588
rect 2280 8576 2286 8628
rect 3050 8576 3056 8628
rect 3108 8616 3114 8628
rect 3145 8619 3203 8625
rect 3145 8616 3157 8619
rect 3108 8588 3157 8616
rect 3108 8576 3114 8588
rect 3145 8585 3157 8588
rect 3191 8585 3203 8619
rect 3145 8579 3203 8585
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5169 8619 5227 8625
rect 5169 8616 5181 8619
rect 5132 8588 5181 8616
rect 5132 8576 5138 8588
rect 5169 8585 5181 8588
rect 5215 8585 5227 8619
rect 5169 8579 5227 8585
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7524 8588 8033 8616
rect 7524 8576 7530 8588
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 10137 8619 10195 8625
rect 10137 8585 10149 8619
rect 10183 8616 10195 8619
rect 10318 8616 10324 8628
rect 10183 8588 10324 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 13078 8616 13084 8628
rect 13039 8588 13084 8616
rect 13078 8576 13084 8588
rect 13136 8576 13142 8628
rect 13170 8576 13176 8628
rect 13228 8616 13234 8628
rect 13265 8619 13323 8625
rect 13265 8616 13277 8619
rect 13228 8588 13277 8616
rect 13228 8576 13234 8588
rect 13265 8585 13277 8588
rect 13311 8585 13323 8619
rect 13446 8616 13452 8628
rect 13407 8588 13452 8616
rect 13265 8579 13323 8585
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 5994 8548 6000 8560
rect 2976 8520 6000 8548
rect 1854 8480 1860 8492
rect 1815 8452 1860 8480
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 2590 8480 2596 8492
rect 2503 8452 2596 8480
rect 2590 8440 2596 8452
rect 2648 8480 2654 8492
rect 2976 8489 3004 8520
rect 5994 8508 6000 8520
rect 6052 8508 6058 8560
rect 6914 8548 6920 8560
rect 6875 8520 6920 8548
rect 6914 8508 6920 8520
rect 6972 8548 6978 8560
rect 9401 8551 9459 8557
rect 6972 8520 9352 8548
rect 6972 8508 6978 8520
rect 2869 8483 2927 8489
rect 2869 8480 2881 8483
rect 2648 8452 2881 8480
rect 2648 8440 2654 8452
rect 2869 8449 2881 8452
rect 2915 8449 2927 8483
rect 2869 8443 2927 8449
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4614 8480 4620 8492
rect 4387 8452 4620 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 1946 8372 1952 8424
rect 2004 8412 2010 8424
rect 2041 8415 2099 8421
rect 2041 8412 2053 8415
rect 2004 8384 2053 8412
rect 2004 8372 2010 8384
rect 2041 8381 2053 8384
rect 2087 8412 2099 8415
rect 2406 8412 2412 8424
rect 2087 8384 2412 8412
rect 2087 8381 2099 8384
rect 2041 8375 2099 8381
rect 2406 8372 2412 8384
rect 2464 8372 2470 8424
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8412 2559 8415
rect 2682 8412 2688 8424
rect 2547 8384 2688 8412
rect 2547 8381 2559 8384
rect 2501 8375 2559 8381
rect 2682 8372 2688 8384
rect 2740 8412 2746 8424
rect 2976 8412 3004 8443
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8449 5503 8483
rect 5445 8443 5503 8449
rect 2740 8384 3004 8412
rect 4249 8415 4307 8421
rect 2740 8372 2746 8384
rect 4249 8381 4261 8415
rect 4295 8412 4307 8415
rect 4295 8384 4568 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 4065 8347 4123 8353
rect 4065 8313 4077 8347
rect 4111 8344 4123 8347
rect 4430 8344 4436 8356
rect 4111 8316 4436 8344
rect 4111 8313 4123 8316
rect 4065 8307 4123 8313
rect 4430 8304 4436 8316
rect 4488 8304 4494 8356
rect 4540 8344 4568 8384
rect 4706 8372 4712 8424
rect 4764 8412 4770 8424
rect 5353 8415 5411 8421
rect 4764 8384 4809 8412
rect 4764 8372 4770 8384
rect 5353 8381 5365 8415
rect 5399 8381 5411 8415
rect 5460 8412 5488 8443
rect 8110 8440 8116 8492
rect 8168 8480 8174 8492
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 8168 8452 8217 8480
rect 8168 8440 8174 8452
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 8205 8443 8263 8449
rect 8312 8452 8493 8480
rect 5718 8412 5724 8424
rect 5460 8384 5724 8412
rect 5353 8375 5411 8381
rect 4724 8344 4752 8372
rect 4540 8316 4752 8344
rect 5368 8344 5396 8375
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 5810 8372 5816 8424
rect 5868 8412 5874 8424
rect 5868 8384 5913 8412
rect 5868 8372 5874 8384
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 8312 8412 8340 8452
rect 8481 8449 8493 8452
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8480 8723 8483
rect 9030 8480 9036 8492
rect 8711 8452 9036 8480
rect 8711 8449 8723 8452
rect 8665 8443 8723 8449
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 9324 8489 9352 8520
rect 9401 8517 9413 8551
rect 9447 8548 9459 8551
rect 11514 8548 11520 8560
rect 9447 8520 11520 8548
rect 9447 8517 9459 8520
rect 9401 8511 9459 8517
rect 11514 8508 11520 8520
rect 11572 8548 11578 8560
rect 11572 8520 11836 8548
rect 11572 8508 11578 8520
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8480 9367 8483
rect 9950 8480 9956 8492
rect 9355 8452 9956 8480
rect 9355 8449 9367 8452
rect 9309 8443 9367 8449
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8480 10379 8483
rect 10502 8480 10508 8492
rect 10367 8452 10508 8480
rect 10367 8449 10379 8452
rect 10321 8443 10379 8449
rect 7432 8384 8340 8412
rect 7432 8372 7438 8384
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 8444 8384 8489 8412
rect 8444 8372 8450 8384
rect 5828 8344 5856 8372
rect 8294 8344 8300 8356
rect 5368 8316 5856 8344
rect 8255 8316 8300 8344
rect 8294 8304 8300 8316
rect 8352 8304 8358 8356
rect 10244 8344 10272 8443
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 11808 8489 11836 8520
rect 12434 8508 12440 8560
rect 12492 8548 12498 8560
rect 13630 8548 13636 8560
rect 12492 8520 13636 8548
rect 12492 8508 12498 8520
rect 13630 8508 13636 8520
rect 13688 8548 13694 8560
rect 14093 8551 14151 8557
rect 14093 8548 14105 8551
rect 13688 8520 14105 8548
rect 13688 8508 13694 8520
rect 14093 8517 14105 8520
rect 14139 8517 14151 8551
rect 14093 8511 14151 8517
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 12618 8440 12624 8492
rect 12676 8480 12682 8492
rect 12894 8480 12900 8492
rect 12676 8452 12900 8480
rect 12676 8440 12682 8452
rect 12894 8440 12900 8452
rect 12952 8480 12958 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 12952 8452 13185 8480
rect 12952 8440 12958 8452
rect 13173 8449 13185 8452
rect 13219 8449 13231 8483
rect 14274 8480 14280 8492
rect 14235 8452 14280 8480
rect 13173 8443 13231 8449
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 15194 8480 15200 8492
rect 15155 8452 15200 8480
rect 15194 8440 15200 8452
rect 15252 8480 15258 8492
rect 15473 8483 15531 8489
rect 15473 8480 15485 8483
rect 15252 8452 15485 8480
rect 15252 8440 15258 8452
rect 15473 8449 15485 8452
rect 15519 8449 15531 8483
rect 15473 8443 15531 8449
rect 12066 8412 12072 8424
rect 12027 8384 12072 8412
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 14461 8415 14519 8421
rect 13320 8384 14136 8412
rect 13320 8372 13326 8384
rect 12897 8347 12955 8353
rect 10244 8316 12434 8344
rect 6454 8236 6460 8288
rect 6512 8276 6518 8288
rect 7009 8279 7067 8285
rect 7009 8276 7021 8279
rect 6512 8248 7021 8276
rect 6512 8236 6518 8248
rect 7009 8245 7021 8248
rect 7055 8245 7067 8279
rect 7009 8239 7067 8245
rect 10505 8279 10563 8285
rect 10505 8245 10517 8279
rect 10551 8276 10563 8279
rect 10870 8276 10876 8288
rect 10551 8248 10876 8276
rect 10551 8245 10563 8248
rect 10505 8239 10563 8245
rect 10870 8236 10876 8248
rect 10928 8236 10934 8288
rect 12406 8276 12434 8316
rect 12897 8313 12909 8347
rect 12943 8344 12955 8347
rect 12986 8344 12992 8356
rect 12943 8316 12992 8344
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 12986 8304 12992 8316
rect 13044 8344 13050 8356
rect 13354 8344 13360 8356
rect 13044 8316 13360 8344
rect 13044 8304 13050 8316
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 14108 8344 14136 8384
rect 14461 8381 14473 8415
rect 14507 8412 14519 8415
rect 15105 8415 15163 8421
rect 15105 8412 15117 8415
rect 14507 8384 15117 8412
rect 14507 8381 14519 8384
rect 14461 8375 14519 8381
rect 15105 8381 15117 8384
rect 15151 8412 15163 8415
rect 15286 8412 15292 8424
rect 15151 8384 15292 8412
rect 15151 8381 15163 8384
rect 15105 8375 15163 8381
rect 15286 8372 15292 8384
rect 15344 8412 15350 8424
rect 15565 8415 15623 8421
rect 15565 8412 15577 8415
rect 15344 8384 15577 8412
rect 15344 8372 15350 8384
rect 15565 8381 15577 8384
rect 15611 8381 15623 8415
rect 15565 8375 15623 8381
rect 14921 8347 14979 8353
rect 14921 8344 14933 8347
rect 14108 8316 14933 8344
rect 14921 8313 14933 8316
rect 14967 8313 14979 8347
rect 14921 8307 14979 8313
rect 12710 8276 12716 8288
rect 12406 8248 12716 8276
rect 12710 8236 12716 8248
rect 12768 8276 12774 8288
rect 13446 8276 13452 8288
rect 12768 8248 13452 8276
rect 12768 8236 12774 8248
rect 13446 8236 13452 8248
rect 13504 8236 13510 8288
rect 1104 8186 16468 8208
rect 1104 8134 3542 8186
rect 3594 8134 3606 8186
rect 3658 8134 3670 8186
rect 3722 8134 3734 8186
rect 3786 8134 8664 8186
rect 8716 8134 8728 8186
rect 8780 8134 8792 8186
rect 8844 8134 8856 8186
rect 8908 8134 13785 8186
rect 13837 8134 13849 8186
rect 13901 8134 13913 8186
rect 13965 8134 13977 8186
rect 14029 8134 16468 8186
rect 1104 8112 16468 8134
rect 2501 8075 2559 8081
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 2590 8072 2596 8084
rect 2547 8044 2596 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 2590 8032 2596 8044
rect 2648 8032 2654 8084
rect 5537 8075 5595 8081
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 6546 8072 6552 8084
rect 5583 8044 6552 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 6641 8075 6699 8081
rect 6641 8041 6653 8075
rect 6687 8072 6699 8075
rect 7374 8072 7380 8084
rect 6687 8044 7380 8072
rect 6687 8041 6699 8044
rect 6641 8035 6699 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 8386 8072 8392 8084
rect 8343 8044 8392 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 10134 8072 10140 8084
rect 9732 8044 10140 8072
rect 9732 8032 9738 8044
rect 10134 8032 10140 8044
rect 10192 8072 10198 8084
rect 12342 8072 12348 8084
rect 10192 8044 10824 8072
rect 12303 8044 12348 8072
rect 10192 8032 10198 8044
rect 6181 8007 6239 8013
rect 6181 7973 6193 8007
rect 6227 8004 6239 8007
rect 8202 8004 8208 8016
rect 6227 7976 8208 8004
rect 6227 7973 6239 7976
rect 6181 7967 6239 7973
rect 8202 7964 8208 7976
rect 8260 7964 8266 8016
rect 9030 8004 9036 8016
rect 8404 7976 9036 8004
rect 4614 7936 4620 7948
rect 4575 7908 4620 7936
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 7374 7936 7380 7948
rect 6012 7908 7380 7936
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7837 2743 7871
rect 2685 7831 2743 7837
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2866 7868 2872 7880
rect 2823 7840 2872 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2700 7800 2728 7831
rect 2866 7828 2872 7840
rect 2924 7868 2930 7880
rect 3053 7871 3111 7877
rect 3053 7868 3065 7871
rect 2924 7840 3065 7868
rect 2924 7828 2930 7840
rect 3053 7837 3065 7840
rect 3099 7868 3111 7871
rect 4157 7871 4215 7877
rect 4157 7868 4169 7871
rect 3099 7840 4169 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 4157 7837 4169 7840
rect 4203 7837 4215 7871
rect 4338 7868 4344 7880
rect 4299 7840 4344 7868
rect 4157 7831 4215 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4430 7828 4436 7880
rect 4488 7868 4494 7880
rect 4488 7840 4533 7868
rect 4488 7828 4494 7840
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 5350 7868 5356 7880
rect 4764 7840 4857 7868
rect 5311 7840 5356 7868
rect 4764 7828 4770 7840
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 6012 7877 6040 7908
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 5997 7871 6055 7877
rect 5997 7837 6009 7871
rect 6043 7837 6055 7871
rect 6638 7868 6644 7880
rect 6599 7840 6644 7868
rect 5997 7831 6055 7837
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7282 7868 7288 7880
rect 6871 7840 7288 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7282 7828 7288 7840
rect 7340 7868 7346 7880
rect 7469 7871 7527 7877
rect 7469 7868 7481 7871
rect 7340 7840 7481 7868
rect 7340 7828 7346 7840
rect 7469 7837 7481 7840
rect 7515 7868 7527 7871
rect 8110 7868 8116 7880
rect 7515 7840 8116 7868
rect 7515 7837 7527 7840
rect 7469 7831 7527 7837
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 8404 7877 8432 7976
rect 9030 7964 9036 7976
rect 9088 8004 9094 8016
rect 10413 8007 10471 8013
rect 10413 8004 10425 8007
rect 9088 7976 10425 8004
rect 9088 7964 9094 7976
rect 10413 7973 10425 7976
rect 10459 7973 10471 8007
rect 10413 7967 10471 7973
rect 10686 7936 10692 7948
rect 9508 7908 10180 7936
rect 10647 7908 10692 7936
rect 9508 7877 9536 7908
rect 10152 7880 10180 7908
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 10796 7945 10824 8044
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 14090 8072 14096 8084
rect 14051 8044 14096 8072
rect 14090 8032 14096 8044
rect 14148 8032 14154 8084
rect 14553 8075 14611 8081
rect 14553 8072 14565 8075
rect 14200 8044 14565 8072
rect 13630 7964 13636 8016
rect 13688 8004 13694 8016
rect 14200 8004 14228 8044
rect 14553 8041 14565 8044
rect 14599 8041 14611 8075
rect 14553 8035 14611 8041
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 15473 8075 15531 8081
rect 15473 8072 15485 8075
rect 15252 8044 15485 8072
rect 15252 8032 15258 8044
rect 15473 8041 15485 8044
rect 15519 8041 15531 8075
rect 15473 8035 15531 8041
rect 15102 8004 15108 8016
rect 13688 7976 14228 8004
rect 14292 7976 15108 8004
rect 13688 7964 13694 7976
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 13354 7936 13360 7948
rect 13035 7908 13360 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7837 9551 7871
rect 9674 7868 9680 7880
rect 9635 7840 9680 7868
rect 9493 7831 9551 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7868 10011 7871
rect 10042 7868 10048 7880
rect 9999 7840 10048 7868
rect 9999 7837 10011 7840
rect 9953 7831 10011 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10134 7828 10140 7880
rect 10192 7868 10198 7880
rect 10597 7871 10655 7877
rect 10597 7868 10609 7871
rect 10192 7840 10609 7868
rect 10192 7828 10198 7840
rect 10597 7837 10609 7840
rect 10643 7837 10655 7871
rect 10597 7831 10655 7837
rect 10870 7828 10876 7880
rect 10928 7868 10934 7880
rect 12437 7871 12495 7877
rect 10928 7840 10973 7868
rect 10928 7828 10934 7840
rect 12437 7837 12449 7871
rect 12483 7868 12495 7871
rect 13078 7868 13084 7880
rect 12483 7840 13084 7868
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 13078 7828 13084 7840
rect 13136 7828 13142 7880
rect 13262 7868 13268 7880
rect 13223 7840 13268 7868
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 14292 7877 14320 7976
rect 15102 7964 15108 7976
rect 15160 7964 15166 8016
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 14366 7828 14372 7880
rect 14424 7868 14430 7880
rect 14642 7868 14648 7880
rect 14424 7840 14469 7868
rect 14603 7840 14648 7868
rect 14424 7828 14430 7840
rect 14642 7828 14648 7840
rect 14700 7828 14706 7880
rect 3145 7803 3203 7809
rect 2700 7772 2774 7800
rect 2746 7744 2774 7772
rect 3145 7769 3157 7803
rect 3191 7769 3203 7803
rect 4724 7800 4752 7828
rect 4724 7772 5672 7800
rect 3145 7763 3203 7769
rect 2746 7704 2780 7744
rect 2774 7692 2780 7704
rect 2832 7732 2838 7744
rect 3160 7732 3188 7763
rect 2832 7704 3188 7732
rect 5644 7732 5672 7772
rect 5810 7760 5816 7812
rect 5868 7800 5874 7812
rect 5868 7772 7420 7800
rect 5868 7760 5874 7772
rect 6730 7732 6736 7744
rect 5644 7704 6736 7732
rect 2832 7692 2838 7704
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 7285 7735 7343 7741
rect 7285 7732 7297 7735
rect 7156 7704 7297 7732
rect 7156 7692 7162 7704
rect 7285 7701 7297 7704
rect 7331 7701 7343 7735
rect 7392 7732 7420 7772
rect 7558 7760 7564 7812
rect 7616 7800 7622 7812
rect 7653 7803 7711 7809
rect 7653 7800 7665 7803
rect 7616 7772 7665 7800
rect 7616 7760 7622 7772
rect 7653 7769 7665 7772
rect 7699 7800 7711 7803
rect 8202 7800 8208 7812
rect 7699 7772 8208 7800
rect 7699 7769 7711 7772
rect 7653 7763 7711 7769
rect 8202 7760 8208 7772
rect 8260 7760 8266 7812
rect 9398 7760 9404 7812
rect 9456 7800 9462 7812
rect 9585 7803 9643 7809
rect 9585 7800 9597 7803
rect 9456 7772 9597 7800
rect 9456 7760 9462 7772
rect 9585 7769 9597 7772
rect 9631 7769 9643 7803
rect 9585 7763 9643 7769
rect 9815 7803 9873 7809
rect 9815 7769 9827 7803
rect 9861 7800 9873 7803
rect 11425 7803 11483 7809
rect 11425 7800 11437 7803
rect 9861 7772 11437 7800
rect 9861 7769 9873 7772
rect 9815 7763 9873 7769
rect 11425 7769 11437 7772
rect 11471 7769 11483 7803
rect 11606 7800 11612 7812
rect 11567 7772 11612 7800
rect 11425 7763 11483 7769
rect 11606 7760 11612 7772
rect 11664 7760 11670 7812
rect 11793 7803 11851 7809
rect 11793 7769 11805 7803
rect 11839 7800 11851 7803
rect 11882 7800 11888 7812
rect 11839 7772 11888 7800
rect 11839 7769 11851 7772
rect 11793 7763 11851 7769
rect 11882 7760 11888 7772
rect 11940 7760 11946 7812
rect 12894 7760 12900 7812
rect 12952 7800 12958 7812
rect 13280 7800 13308 7828
rect 12952 7772 13308 7800
rect 13541 7803 13599 7809
rect 12952 7760 12958 7772
rect 13541 7769 13553 7803
rect 13587 7800 13599 7803
rect 14826 7800 14832 7812
rect 13587 7772 14832 7800
rect 13587 7769 13599 7772
rect 13541 7763 13599 7769
rect 14826 7760 14832 7772
rect 14884 7800 14890 7812
rect 15105 7803 15163 7809
rect 15105 7800 15117 7803
rect 14884 7772 15117 7800
rect 14884 7760 14890 7772
rect 15105 7769 15117 7772
rect 15151 7769 15163 7803
rect 15286 7800 15292 7812
rect 15247 7772 15292 7800
rect 15105 7763 15163 7769
rect 15286 7760 15292 7772
rect 15344 7760 15350 7812
rect 9309 7735 9367 7741
rect 9309 7732 9321 7735
rect 7392 7704 9321 7732
rect 7285 7695 7343 7701
rect 9309 7701 9321 7704
rect 9355 7701 9367 7735
rect 9309 7695 9367 7701
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 12434 7732 12440 7744
rect 10652 7704 12440 7732
rect 10652 7692 10658 7704
rect 12434 7692 12440 7704
rect 12492 7692 12498 7744
rect 13078 7692 13084 7744
rect 13136 7732 13142 7744
rect 13173 7735 13231 7741
rect 13173 7732 13185 7735
rect 13136 7704 13185 7732
rect 13136 7692 13142 7704
rect 13173 7701 13185 7704
rect 13219 7701 13231 7735
rect 13173 7695 13231 7701
rect 13357 7735 13415 7741
rect 13357 7701 13369 7735
rect 13403 7732 13415 7735
rect 13446 7732 13452 7744
rect 13403 7704 13452 7732
rect 13403 7701 13415 7704
rect 13357 7695 13415 7701
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 1104 7642 16468 7664
rect 1104 7590 6103 7642
rect 6155 7590 6167 7642
rect 6219 7590 6231 7642
rect 6283 7590 6295 7642
rect 6347 7590 11224 7642
rect 11276 7590 11288 7642
rect 11340 7590 11352 7642
rect 11404 7590 11416 7642
rect 11468 7590 16468 7642
rect 1104 7568 16468 7590
rect 1854 7488 1860 7540
rect 1912 7528 1918 7540
rect 2225 7531 2283 7537
rect 2225 7528 2237 7531
rect 1912 7500 2237 7528
rect 1912 7488 1918 7500
rect 2225 7497 2237 7500
rect 2271 7497 2283 7531
rect 2225 7491 2283 7497
rect 4157 7531 4215 7537
rect 4157 7497 4169 7531
rect 4203 7497 4215 7531
rect 4157 7491 4215 7497
rect 2682 7460 2688 7472
rect 2424 7432 2688 7460
rect 2424 7401 2452 7432
rect 2682 7420 2688 7432
rect 2740 7420 2746 7472
rect 4172 7460 4200 7491
rect 4614 7488 4620 7540
rect 4672 7528 4678 7540
rect 5261 7531 5319 7537
rect 5261 7528 5273 7531
rect 4672 7500 5273 7528
rect 4672 7488 4678 7500
rect 5261 7497 5273 7500
rect 5307 7497 5319 7531
rect 6914 7528 6920 7540
rect 5261 7491 5319 7497
rect 5368 7500 6920 7528
rect 5368 7460 5396 7500
rect 6914 7488 6920 7500
rect 6972 7488 6978 7540
rect 7466 7528 7472 7540
rect 7024 7500 7472 7528
rect 7024 7469 7052 7500
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 7852 7500 8236 7528
rect 7009 7463 7067 7469
rect 7009 7460 7021 7463
rect 4172 7432 5396 7460
rect 6564 7432 7021 7460
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7361 2467 7395
rect 2409 7355 2467 7361
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 2590 7392 2596 7404
rect 2547 7364 2596 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2590 7352 2596 7364
rect 2648 7352 2654 7404
rect 2774 7352 2780 7404
rect 2832 7392 2838 7404
rect 3970 7392 3976 7404
rect 2832 7364 2877 7392
rect 3931 7364 3976 7392
rect 2832 7352 2838 7364
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 4614 7392 4620 7404
rect 4575 7364 4620 7392
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 6564 7401 6592 7432
rect 7009 7429 7021 7432
rect 7055 7429 7067 7463
rect 7742 7460 7748 7472
rect 7703 7432 7748 7460
rect 7009 7423 7067 7429
rect 7742 7420 7748 7432
rect 7800 7420 7806 7472
rect 7852 7469 7880 7500
rect 7837 7463 7895 7469
rect 7837 7429 7849 7463
rect 7883 7429 7895 7463
rect 8208 7460 8236 7500
rect 8386 7488 8392 7540
rect 8444 7528 8450 7540
rect 8757 7531 8815 7537
rect 8757 7528 8769 7531
rect 8444 7500 8769 7528
rect 8444 7488 8450 7500
rect 8757 7497 8769 7500
rect 8803 7497 8815 7531
rect 9674 7528 9680 7540
rect 8757 7491 8815 7497
rect 8864 7500 9680 7528
rect 8864 7460 8892 7500
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7528 10011 7531
rect 10134 7528 10140 7540
rect 9999 7500 10140 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 12158 7528 12164 7540
rect 11716 7500 12164 7528
rect 10594 7460 10600 7472
rect 8208 7432 8892 7460
rect 9416 7432 10600 7460
rect 7837 7423 7895 7429
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 5859 7364 6561 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7324 2743 7327
rect 2866 7324 2872 7336
rect 2731 7296 2872 7324
rect 2731 7293 2743 7296
rect 2685 7287 2743 7293
rect 2866 7284 2872 7296
rect 2924 7284 2930 7336
rect 4798 7256 4804 7268
rect 4759 7228 4804 7256
rect 4798 7216 4804 7228
rect 4856 7216 4862 7268
rect 5460 7256 5488 7355
rect 5552 7324 5580 7355
rect 5718 7324 5724 7336
rect 5552 7296 5724 7324
rect 5718 7284 5724 7296
rect 5776 7324 5782 7336
rect 6656 7324 6684 7355
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 7466 7392 7472 7404
rect 6788 7364 7472 7392
rect 6788 7352 6794 7364
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 7650 7392 7656 7404
rect 7611 7364 7656 7392
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 7926 7352 7932 7404
rect 7984 7401 7990 7404
rect 7984 7395 8033 7401
rect 7984 7361 7987 7395
rect 8021 7361 8033 7395
rect 7984 7355 8033 7361
rect 7984 7352 7990 7355
rect 8478 7352 8484 7404
rect 8536 7392 8542 7404
rect 9416 7401 9444 7432
rect 10594 7420 10600 7432
rect 10652 7420 10658 7472
rect 10689 7463 10747 7469
rect 10689 7429 10701 7463
rect 10735 7460 10747 7463
rect 11517 7463 11575 7469
rect 11517 7460 11529 7463
rect 10735 7432 11529 7460
rect 10735 7429 10747 7432
rect 10689 7423 10747 7429
rect 11517 7429 11529 7432
rect 11563 7429 11575 7463
rect 11517 7423 11575 7429
rect 8573 7395 8631 7401
rect 8573 7392 8585 7395
rect 8536 7364 8585 7392
rect 8536 7352 8542 7364
rect 8573 7361 8585 7364
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7361 9459 7395
rect 10042 7392 10048 7404
rect 10003 7364 10048 7392
rect 9401 7355 9459 7361
rect 10042 7352 10048 7364
rect 10100 7392 10106 7404
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 10100 7364 10517 7392
rect 10100 7352 10106 7364
rect 10505 7361 10517 7364
rect 10551 7361 10563 7395
rect 10870 7392 10876 7404
rect 10831 7364 10876 7392
rect 10505 7355 10563 7361
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 10962 7352 10968 7404
rect 11020 7392 11026 7404
rect 11716 7401 11744 7500
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 13814 7488 13820 7540
rect 13872 7528 13878 7540
rect 14090 7528 14096 7540
rect 13872 7500 14096 7528
rect 13872 7488 13878 7500
rect 14090 7488 14096 7500
rect 14148 7528 14154 7540
rect 14734 7528 14740 7540
rect 14148 7500 14740 7528
rect 14148 7488 14154 7500
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 15105 7531 15163 7537
rect 15105 7497 15117 7531
rect 15151 7528 15163 7531
rect 15286 7528 15292 7540
rect 15151 7500 15292 7528
rect 15151 7497 15163 7500
rect 15105 7491 15163 7497
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 13170 7460 13176 7472
rect 12084 7432 13176 7460
rect 12084 7404 12112 7432
rect 13170 7420 13176 7432
rect 13228 7420 13234 7472
rect 14752 7460 14780 7488
rect 14752 7432 15608 7460
rect 11701 7395 11759 7401
rect 11020 7364 11652 7392
rect 11020 7352 11026 7364
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 5776 7296 6408 7324
rect 5776 7284 5782 7296
rect 5810 7256 5816 7268
rect 5460 7228 5816 7256
rect 5810 7216 5816 7228
rect 5868 7216 5874 7268
rect 6380 7265 6408 7296
rect 6656 7296 6929 7324
rect 6365 7259 6423 7265
rect 6365 7225 6377 7259
rect 6411 7225 6423 7259
rect 6365 7219 6423 7225
rect 5721 7191 5779 7197
rect 5721 7157 5733 7191
rect 5767 7188 5779 7191
rect 6656 7188 6684 7296
rect 6917 7293 6929 7296
rect 6963 7324 6975 7327
rect 7006 7324 7012 7336
rect 6963 7296 7012 7324
rect 6963 7293 6975 7296
rect 6917 7287 6975 7293
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 8113 7327 8171 7333
rect 8113 7324 8125 7327
rect 8036 7296 8125 7324
rect 7098 7216 7104 7268
rect 7156 7256 7162 7268
rect 7156 7228 7880 7256
rect 7156 7216 7162 7228
rect 7466 7188 7472 7200
rect 5767 7160 6684 7188
rect 7427 7160 7472 7188
rect 5767 7157 5779 7160
rect 5721 7151 5779 7157
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 7852 7188 7880 7228
rect 8036 7188 8064 7296
rect 8113 7293 8125 7296
rect 8159 7293 8171 7327
rect 8113 7287 8171 7293
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 11054 7324 11060 7336
rect 8352 7296 11060 7324
rect 8352 7284 8358 7296
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 11624 7324 11652 7364
rect 11701 7361 11713 7395
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7392 11851 7395
rect 11974 7392 11980 7404
rect 11839 7364 11980 7392
rect 11839 7361 11851 7364
rect 11793 7355 11851 7361
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12124 7364 12217 7392
rect 12124 7352 12130 7364
rect 12250 7352 12256 7404
rect 12308 7392 12314 7404
rect 12529 7395 12587 7401
rect 12529 7392 12541 7395
rect 12308 7364 12541 7392
rect 12308 7352 12314 7364
rect 12529 7361 12541 7364
rect 12575 7361 12587 7395
rect 12710 7392 12716 7404
rect 12671 7364 12716 7392
rect 12529 7355 12587 7361
rect 12710 7352 12716 7364
rect 12768 7352 12774 7404
rect 13814 7392 13820 7404
rect 13775 7364 13820 7392
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 14550 7392 14556 7404
rect 14511 7364 14556 7392
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 14734 7352 14740 7404
rect 14792 7392 14798 7404
rect 14829 7395 14887 7401
rect 14829 7392 14841 7395
rect 14792 7364 14841 7392
rect 14792 7352 14798 7364
rect 14829 7361 14841 7364
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 14921 7395 14979 7401
rect 14921 7361 14933 7395
rect 14967 7392 14979 7395
rect 15102 7392 15108 7404
rect 14967 7364 15108 7392
rect 14967 7361 14979 7364
rect 14921 7355 14979 7361
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 15580 7401 15608 7432
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7361 15623 7395
rect 15565 7355 15623 7361
rect 12084 7324 12112 7352
rect 12618 7324 12624 7336
rect 11624 7296 12112 7324
rect 12406 7296 12624 7324
rect 9030 7216 9036 7268
rect 9088 7256 9094 7268
rect 12406 7256 12434 7296
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 14366 7284 14372 7336
rect 14424 7324 14430 7336
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 14424 7296 14657 7324
rect 14424 7284 14430 7296
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 14645 7287 14703 7293
rect 9088 7228 12434 7256
rect 9088 7216 9094 7228
rect 7852 7160 8064 7188
rect 8110 7148 8116 7200
rect 8168 7188 8174 7200
rect 9217 7191 9275 7197
rect 9217 7188 9229 7191
rect 8168 7160 9229 7188
rect 8168 7148 8174 7160
rect 9217 7157 9229 7160
rect 9263 7188 9275 7191
rect 11606 7188 11612 7200
rect 9263 7160 11612 7188
rect 9263 7157 9275 7160
rect 9217 7151 9275 7157
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 11977 7191 12035 7197
rect 11977 7188 11989 7191
rect 11756 7160 11989 7188
rect 11756 7148 11762 7160
rect 11977 7157 11989 7160
rect 12023 7157 12035 7191
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 11977 7151 12035 7157
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13354 7148 13360 7200
rect 13412 7188 13418 7200
rect 13633 7191 13691 7197
rect 13633 7188 13645 7191
rect 13412 7160 13645 7188
rect 13412 7148 13418 7160
rect 13633 7157 13645 7160
rect 13679 7157 13691 7191
rect 13633 7151 13691 7157
rect 14550 7148 14556 7200
rect 14608 7188 14614 7200
rect 15657 7191 15715 7197
rect 15657 7188 15669 7191
rect 14608 7160 15669 7188
rect 14608 7148 14614 7160
rect 15657 7157 15669 7160
rect 15703 7157 15715 7191
rect 15657 7151 15715 7157
rect 1104 7098 16468 7120
rect 1104 7046 3542 7098
rect 3594 7046 3606 7098
rect 3658 7046 3670 7098
rect 3722 7046 3734 7098
rect 3786 7046 8664 7098
rect 8716 7046 8728 7098
rect 8780 7046 8792 7098
rect 8844 7046 8856 7098
rect 8908 7046 13785 7098
rect 13837 7046 13849 7098
rect 13901 7046 13913 7098
rect 13965 7046 13977 7098
rect 14029 7046 16468 7098
rect 1104 7024 16468 7046
rect 2406 6984 2412 6996
rect 2367 6956 2412 6984
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 2774 6944 2780 6996
rect 2832 6984 2838 6996
rect 3789 6987 3847 6993
rect 3789 6984 3801 6987
rect 2832 6956 3801 6984
rect 2832 6944 2838 6956
rect 3789 6953 3801 6956
rect 3835 6953 3847 6987
rect 7466 6984 7472 6996
rect 3789 6947 3847 6953
rect 6288 6956 7472 6984
rect 6288 6916 6316 6956
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 7616 6956 10824 6984
rect 7616 6944 7622 6956
rect 8018 6916 8024 6928
rect 6012 6888 6316 6916
rect 6932 6888 7328 6916
rect 7979 6888 8024 6916
rect 2593 6851 2651 6857
rect 2593 6817 2605 6851
rect 2639 6848 2651 6851
rect 3973 6851 4031 6857
rect 2639 6820 3372 6848
rect 2639 6817 2651 6820
rect 2593 6811 2651 6817
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6780 1455 6783
rect 2685 6783 2743 6789
rect 1443 6752 2452 6780
rect 1443 6749 1455 6752
rect 1397 6743 1455 6749
rect 2424 6712 2452 6752
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2731 6752 2973 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 2961 6749 2973 6752
rect 3007 6780 3019 6783
rect 3234 6780 3240 6792
rect 3007 6752 3240 6780
rect 3007 6749 3019 6752
rect 2961 6743 3019 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 2866 6712 2872 6724
rect 2424 6684 2872 6712
rect 2866 6672 2872 6684
rect 2924 6672 2930 6724
rect 3050 6672 3056 6724
rect 3108 6712 3114 6724
rect 3344 6712 3372 6820
rect 3973 6817 3985 6851
rect 4019 6848 4031 6851
rect 4433 6851 4491 6857
rect 4433 6848 4445 6851
rect 4019 6820 4445 6848
rect 4019 6817 4031 6820
rect 3973 6811 4031 6817
rect 4433 6817 4445 6820
rect 4479 6848 4491 6851
rect 4522 6848 4528 6860
rect 4479 6820 4528 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 4522 6808 4528 6820
rect 4580 6848 4586 6860
rect 6012 6848 6040 6888
rect 4580 6820 6040 6848
rect 6089 6851 6147 6857
rect 4580 6808 4586 6820
rect 6089 6817 6101 6851
rect 6135 6848 6147 6851
rect 6932 6848 6960 6888
rect 7098 6848 7104 6860
rect 6135 6820 6960 6848
rect 7059 6820 7104 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6780 4123 6783
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 4111 6752 4353 6780
rect 4111 6749 4123 6752
rect 4065 6743 4123 6749
rect 4341 6749 4353 6752
rect 4387 6780 4399 6783
rect 4890 6780 4896 6792
rect 4387 6752 4896 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 5442 6780 5448 6792
rect 5399 6752 5448 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6780 5595 6783
rect 5902 6780 5908 6792
rect 5583 6752 5908 6780
rect 5583 6749 5595 6752
rect 5537 6743 5595 6749
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 6638 6780 6644 6792
rect 6227 6752 6644 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 6822 6780 6828 6792
rect 6783 6752 6828 6780
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 7300 6789 7328 6888
rect 8018 6876 8024 6888
rect 8076 6876 8082 6928
rect 10686 6916 10692 6928
rect 10152 6888 10692 6916
rect 8113 6851 8171 6857
rect 8113 6848 8125 6851
rect 7852 6820 8125 6848
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 7285 6783 7343 6789
rect 7055 6749 7072 6780
rect 7009 6743 7072 6749
rect 7285 6749 7297 6783
rect 7331 6780 7343 6783
rect 7466 6780 7472 6792
rect 7331 6752 7472 6780
rect 7331 6749 7343 6752
rect 7285 6743 7343 6749
rect 3108 6684 6132 6712
rect 3108 6672 3114 6684
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 1670 6604 1676 6656
rect 1728 6644 1734 6656
rect 5350 6644 5356 6656
rect 1728 6616 5356 6644
rect 1728 6604 1734 6616
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 5442 6604 5448 6656
rect 5500 6644 5506 6656
rect 6104 6644 6132 6684
rect 6641 6647 6699 6653
rect 6641 6644 6653 6647
rect 5500 6616 5545 6644
rect 6104 6616 6653 6644
rect 5500 6604 5506 6616
rect 6641 6613 6653 6616
rect 6687 6613 6699 6647
rect 6932 6644 6960 6743
rect 7044 6712 7072 6743
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 7852 6712 7880 6820
rect 8113 6817 8125 6820
rect 8159 6848 8171 6851
rect 8754 6848 8760 6860
rect 8159 6820 8760 6848
rect 8159 6817 8171 6820
rect 8113 6811 8171 6817
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 9999 6851 10057 6857
rect 9456 6820 9674 6848
rect 9456 6808 9462 6820
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 7044 6684 7880 6712
rect 7282 6644 7288 6656
rect 6932 6616 7288 6644
rect 6641 6607 6699 6613
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 7650 6604 7656 6656
rect 7708 6644 7714 6656
rect 7745 6647 7803 6653
rect 7745 6644 7757 6647
rect 7708 6616 7757 6644
rect 7708 6604 7714 6616
rect 7745 6613 7757 6616
rect 7791 6613 7803 6647
rect 7944 6644 7972 6743
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 8260 6752 8305 6780
rect 8260 6740 8266 6752
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 9493 6783 9551 6789
rect 8444 6752 8489 6780
rect 8444 6740 8450 6752
rect 9493 6749 9505 6783
rect 9539 6749 9551 6783
rect 9646 6780 9674 6820
rect 9999 6817 10011 6851
rect 10045 6848 10057 6851
rect 10152 6848 10180 6888
rect 10686 6876 10692 6888
rect 10744 6876 10750 6928
rect 10796 6916 10824 6956
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 12066 6984 12072 6996
rect 11112 6956 12072 6984
rect 11112 6944 11118 6956
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 12805 6987 12863 6993
rect 12805 6984 12817 6987
rect 12176 6956 12817 6984
rect 12176 6916 12204 6956
rect 12805 6953 12817 6956
rect 12851 6953 12863 6987
rect 12805 6947 12863 6953
rect 10796 6888 12204 6916
rect 13170 6876 13176 6928
rect 13228 6916 13234 6928
rect 13228 6888 13676 6916
rect 13228 6876 13234 6888
rect 10045 6820 10180 6848
rect 10045 6817 10057 6820
rect 9999 6811 10057 6817
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 11333 6851 11391 6857
rect 11333 6848 11345 6851
rect 10376 6820 11345 6848
rect 10376 6808 10382 6820
rect 11333 6817 11345 6820
rect 11379 6817 11391 6851
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 11333 6811 11391 6817
rect 13004 6820 13461 6848
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 9646 6779 9904 6780
rect 10152 6779 10241 6780
rect 9646 6752 10241 6779
rect 9876 6751 10180 6752
rect 9493 6743 9551 6749
rect 10229 6749 10241 6752
rect 10275 6780 10287 6783
rect 11701 6783 11759 6789
rect 11701 6782 11713 6783
rect 11440 6780 11560 6782
rect 10275 6752 11008 6780
rect 10275 6749 10287 6752
rect 10229 6743 10287 6749
rect 9508 6712 9536 6743
rect 10870 6712 10876 6724
rect 9508 6684 10876 6712
rect 10870 6672 10876 6684
rect 10928 6672 10934 6724
rect 10980 6712 11008 6752
rect 11348 6779 11560 6780
rect 11624 6779 11713 6782
rect 11348 6754 11713 6779
rect 11348 6752 11468 6754
rect 11348 6712 11376 6752
rect 11532 6751 11652 6754
rect 11701 6749 11713 6754
rect 11747 6749 11759 6783
rect 11701 6743 11759 6749
rect 11790 6740 11796 6792
rect 11848 6780 11854 6792
rect 13004 6789 13032 6820
rect 13449 6817 13461 6820
rect 13495 6848 13507 6851
rect 13538 6848 13544 6860
rect 13495 6820 13544 6848
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 11977 6783 12035 6789
rect 11848 6752 11893 6780
rect 11848 6740 11854 6752
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 12989 6783 13047 6789
rect 12989 6780 13001 6783
rect 12023 6752 13001 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12989 6749 13001 6752
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6780 13139 6783
rect 13648 6780 13676 6888
rect 14366 6848 14372 6860
rect 14200 6820 14372 6848
rect 14200 6789 14228 6820
rect 14366 6808 14372 6820
rect 14424 6808 14430 6860
rect 15378 6848 15384 6860
rect 15212 6820 15384 6848
rect 15212 6789 15240 6820
rect 15378 6808 15384 6820
rect 15436 6848 15442 6860
rect 15657 6851 15715 6857
rect 15657 6848 15669 6851
rect 15436 6820 15669 6848
rect 15436 6808 15442 6820
rect 15657 6817 15669 6820
rect 15703 6817 15715 6851
rect 15657 6811 15715 6817
rect 14185 6783 14243 6789
rect 14185 6780 14197 6783
rect 13127 6752 13216 6780
rect 13648 6752 14197 6780
rect 13127 6749 13139 6752
rect 13081 6743 13139 6749
rect 13188 6724 13216 6752
rect 14185 6749 14197 6752
rect 14231 6749 14243 6783
rect 14185 6743 14243 6749
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 15197 6783 15255 6789
rect 15197 6780 15209 6783
rect 14599 6752 15209 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 15197 6749 15209 6752
rect 15243 6749 15255 6783
rect 15197 6743 15255 6749
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 15565 6783 15623 6789
rect 15565 6780 15577 6783
rect 15344 6752 15577 6780
rect 15344 6740 15350 6752
rect 15565 6749 15577 6752
rect 15611 6749 15623 6783
rect 15565 6743 15623 6749
rect 10980 6684 11376 6712
rect 11422 6672 11428 6724
rect 11480 6721 11486 6724
rect 11480 6715 11529 6721
rect 11480 6681 11483 6715
rect 11517 6681 11529 6715
rect 11480 6675 11529 6681
rect 11596 6715 11654 6721
rect 11596 6681 11608 6715
rect 11642 6712 11654 6715
rect 11642 6684 11836 6712
rect 11642 6681 11654 6684
rect 11596 6675 11654 6681
rect 11480 6672 11486 6675
rect 11808 6656 11836 6684
rect 13170 6672 13176 6724
rect 13228 6712 13234 6724
rect 13357 6715 13415 6721
rect 13357 6712 13369 6715
rect 13228 6684 13369 6712
rect 13228 6672 13234 6684
rect 13357 6681 13369 6684
rect 13403 6681 13415 6715
rect 13357 6675 13415 6681
rect 14274 6672 14280 6724
rect 14332 6712 14338 6724
rect 14369 6715 14427 6721
rect 14369 6712 14381 6715
rect 14332 6684 14381 6712
rect 14332 6672 14338 6684
rect 14369 6681 14381 6684
rect 14415 6681 14427 6715
rect 14369 6675 14427 6681
rect 8018 6644 8024 6656
rect 7931 6616 8024 6644
rect 7745 6607 7803 6613
rect 8018 6604 8024 6616
rect 8076 6644 8082 6656
rect 9309 6647 9367 6653
rect 9309 6644 9321 6647
rect 8076 6616 9321 6644
rect 8076 6604 8082 6616
rect 9309 6613 9321 6616
rect 9355 6644 9367 6647
rect 10962 6644 10968 6656
rect 9355 6616 10968 6644
rect 9355 6613 9367 6616
rect 9309 6607 9367 6613
rect 10962 6604 10968 6616
rect 11020 6604 11026 6656
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 13078 6644 13084 6656
rect 11848 6616 13084 6644
rect 11848 6604 11854 6616
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 15010 6644 15016 6656
rect 14971 6616 15016 6644
rect 15010 6604 15016 6616
rect 15068 6604 15074 6656
rect 1104 6554 16468 6576
rect 1104 6502 6103 6554
rect 6155 6502 6167 6554
rect 6219 6502 6231 6554
rect 6283 6502 6295 6554
rect 6347 6502 11224 6554
rect 11276 6502 11288 6554
rect 11340 6502 11352 6554
rect 11404 6502 11416 6554
rect 11468 6502 16468 6554
rect 1104 6480 16468 6502
rect 3234 6440 3240 6452
rect 3195 6412 3240 6440
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 4890 6440 4896 6452
rect 3344 6412 4016 6440
rect 4851 6412 4896 6440
rect 1578 6332 1584 6384
rect 1636 6372 1642 6384
rect 3344 6372 3372 6412
rect 3988 6372 4016 6412
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 5442 6400 5448 6452
rect 5500 6440 5506 6452
rect 7926 6440 7932 6452
rect 5500 6412 7932 6440
rect 5500 6400 5506 6412
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 8113 6443 8171 6449
rect 8113 6409 8125 6443
rect 8159 6440 8171 6443
rect 8202 6440 8208 6452
rect 8159 6412 8208 6440
rect 8159 6409 8171 6412
rect 8113 6403 8171 6409
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 8754 6440 8760 6452
rect 8715 6412 8760 6440
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 12066 6440 12072 6452
rect 8864 6412 11928 6440
rect 12027 6412 12072 6440
rect 8864 6372 8892 6412
rect 1636 6344 3372 6372
rect 3436 6344 3924 6372
rect 3988 6344 8892 6372
rect 9401 6375 9459 6381
rect 1636 6332 1642 6344
rect 1670 6304 1676 6316
rect 1631 6276 1676 6304
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 3436 6313 3464 6344
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 3528 6236 3556 6267
rect 3786 6236 3792 6248
rect 3528 6208 3792 6236
rect 3786 6196 3792 6208
rect 3844 6196 3850 6248
rect 3896 6245 3924 6344
rect 9401 6341 9413 6375
rect 9447 6372 9459 6375
rect 9674 6372 9680 6384
rect 9447 6344 9680 6372
rect 9447 6341 9459 6344
rect 9401 6335 9459 6341
rect 9674 6332 9680 6344
rect 9732 6372 9738 6384
rect 10686 6372 10692 6384
rect 9732 6344 10088 6372
rect 9732 6332 9738 6344
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6304 4859 6307
rect 5169 6307 5227 6313
rect 5169 6304 5181 6307
rect 4847 6276 5181 6304
rect 4847 6273 4859 6276
rect 4801 6267 4859 6273
rect 5169 6273 5181 6276
rect 5215 6273 5227 6307
rect 6546 6304 6552 6316
rect 5169 6267 5227 6273
rect 5276 6276 5580 6304
rect 6507 6276 6552 6304
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4430 6236 4436 6248
rect 3927 6208 4436 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6236 5135 6239
rect 5276 6236 5304 6276
rect 5552 6248 5580 6276
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 6880 6276 7205 6304
rect 6880 6264 6886 6276
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6304 7435 6307
rect 7834 6304 7840 6316
rect 7423 6276 7840 6304
rect 7423 6273 7435 6276
rect 7377 6267 7435 6273
rect 5442 6236 5448 6248
rect 5123 6208 5304 6236
rect 5403 6208 5448 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 5534 6196 5540 6248
rect 5592 6236 5598 6248
rect 6457 6239 6515 6245
rect 5592 6208 5637 6236
rect 5592 6196 5598 6208
rect 6457 6205 6469 6239
rect 6503 6236 6515 6239
rect 6638 6236 6644 6248
rect 6503 6208 6644 6236
rect 6503 6205 6515 6208
rect 6457 6199 6515 6205
rect 6638 6196 6644 6208
rect 6696 6196 6702 6248
rect 7006 6236 7012 6248
rect 6967 6208 7012 6236
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 7208 6236 7236 6267
rect 7834 6264 7840 6276
rect 7892 6264 7898 6316
rect 8018 6304 8024 6316
rect 7979 6276 8024 6304
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 8036 6236 8064 6264
rect 7208 6208 8064 6236
rect 8220 6236 8248 6267
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8444 6276 8861 6304
rect 8444 6264 8450 6276
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6304 9551 6307
rect 9766 6304 9772 6316
rect 9539 6276 9772 6304
rect 9539 6273 9551 6276
rect 9493 6267 9551 6273
rect 8294 6236 8300 6248
rect 8220 6208 8300 6236
rect 8294 6196 8300 6208
rect 8352 6236 8358 6248
rect 8478 6236 8484 6248
rect 8352 6208 8484 6236
rect 8352 6196 8358 6208
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 8864 6236 8892 6267
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 8864 6208 9965 6236
rect 9953 6205 9965 6208
rect 9999 6205 10011 6239
rect 10060 6236 10088 6344
rect 10336 6344 10692 6372
rect 10336 6326 10364 6344
rect 10686 6332 10692 6344
rect 10744 6372 10750 6384
rect 11422 6372 11428 6384
rect 10744 6344 11428 6372
rect 10744 6332 10750 6344
rect 11422 6332 11428 6344
rect 11480 6332 11486 6384
rect 10244 6313 10364 6326
rect 10229 6307 10364 6313
rect 10229 6273 10241 6307
rect 10275 6298 10364 6307
rect 10413 6310 10471 6313
rect 10413 6307 10548 6310
rect 10275 6273 10287 6298
rect 10229 6267 10287 6273
rect 10413 6273 10425 6307
rect 10459 6304 10548 6307
rect 10778 6304 10784 6316
rect 10459 6282 10784 6304
rect 10459 6273 10471 6282
rect 10520 6276 10784 6282
rect 10413 6267 10471 6273
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 11900 6304 11928 6412
rect 12066 6400 12072 6412
rect 12124 6400 12130 6452
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 14642 6440 14648 6452
rect 12216 6412 14648 6440
rect 12216 6400 12222 6412
rect 14642 6400 14648 6412
rect 14700 6400 14706 6452
rect 12253 6375 12311 6381
rect 12253 6341 12265 6375
rect 12299 6372 12311 6375
rect 12894 6372 12900 6384
rect 12299 6344 12900 6372
rect 12299 6341 12311 6344
rect 12253 6335 12311 6341
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 14458 6332 14464 6384
rect 14516 6372 14522 6384
rect 14737 6375 14795 6381
rect 14737 6372 14749 6375
rect 14516 6344 14749 6372
rect 14516 6332 14522 6344
rect 14737 6341 14749 6344
rect 14783 6341 14795 6375
rect 14737 6335 14795 6341
rect 12342 6304 12348 6316
rect 11900 6276 12348 6304
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12802 6304 12808 6316
rect 12483 6276 12808 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 12802 6264 12808 6276
rect 12860 6304 12866 6316
rect 13081 6307 13139 6313
rect 13081 6304 13093 6307
rect 12860 6276 13093 6304
rect 12860 6264 12866 6276
rect 13081 6273 13093 6276
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 13357 6307 13415 6313
rect 13357 6304 13369 6307
rect 13228 6276 13369 6304
rect 13228 6264 13234 6276
rect 13357 6273 13369 6276
rect 13403 6273 13415 6307
rect 13538 6304 13544 6316
rect 13499 6276 13544 6304
rect 13357 6267 13415 6273
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 13722 6264 13728 6316
rect 13780 6304 13786 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 13780 6276 14105 6304
rect 13780 6264 13786 6276
rect 14093 6273 14105 6276
rect 14139 6273 14151 6307
rect 14918 6304 14924 6316
rect 14879 6276 14924 6304
rect 14093 6267 14151 6273
rect 14918 6264 14924 6276
rect 14976 6264 14982 6316
rect 15197 6307 15255 6313
rect 15197 6273 15209 6307
rect 15243 6273 15255 6307
rect 15378 6304 15384 6316
rect 15339 6276 15384 6304
rect 15197 6267 15255 6273
rect 10137 6239 10195 6245
rect 10137 6236 10149 6239
rect 10060 6208 10149 6236
rect 9953 6199 10011 6205
rect 10137 6205 10149 6208
rect 10183 6205 10195 6239
rect 10137 6199 10195 6205
rect 10318 6196 10324 6248
rect 10376 6236 10382 6248
rect 15212 6236 15240 6267
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 15286 6236 15292 6248
rect 10376 6208 10421 6236
rect 15212 6208 15292 6236
rect 10376 6196 10382 6208
rect 15286 6196 15292 6208
rect 15344 6196 15350 6248
rect 2774 6128 2780 6180
rect 2832 6168 2838 6180
rect 9766 6168 9772 6180
rect 2832 6140 9772 6168
rect 2832 6128 2838 6140
rect 9766 6128 9772 6140
rect 9824 6128 9830 6180
rect 14274 6168 14280 6180
rect 14235 6140 14280 6168
rect 14274 6128 14280 6140
rect 14332 6128 14338 6180
rect 4801 6103 4859 6109
rect 4801 6069 4813 6103
rect 4847 6100 4859 6103
rect 5442 6100 5448 6112
rect 4847 6072 5448 6100
rect 4847 6069 4859 6072
rect 4801 6063 4859 6069
rect 5442 6060 5448 6072
rect 5500 6100 5506 6112
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 5500 6072 12909 6100
rect 5500 6060 5506 6072
rect 12897 6069 12909 6072
rect 12943 6069 12955 6103
rect 12897 6063 12955 6069
rect 1104 6010 16468 6032
rect 1104 5958 3542 6010
rect 3594 5958 3606 6010
rect 3658 5958 3670 6010
rect 3722 5958 3734 6010
rect 3786 5958 8664 6010
rect 8716 5958 8728 6010
rect 8780 5958 8792 6010
rect 8844 5958 8856 6010
rect 8908 5958 13785 6010
rect 13837 5958 13849 6010
rect 13901 5958 13913 6010
rect 13965 5958 13977 6010
rect 14029 5958 16468 6010
rect 1104 5936 16468 5958
rect 3145 5899 3203 5905
rect 3145 5865 3157 5899
rect 3191 5896 3203 5899
rect 3878 5896 3884 5908
rect 3191 5868 3884 5896
rect 3191 5865 3203 5868
rect 3145 5859 3203 5865
rect 3878 5856 3884 5868
rect 3936 5896 3942 5908
rect 4341 5899 4399 5905
rect 4341 5896 4353 5899
rect 3936 5868 4353 5896
rect 3936 5856 3942 5868
rect 4341 5865 4353 5868
rect 4387 5865 4399 5899
rect 4341 5859 4399 5865
rect 4430 5856 4436 5908
rect 4488 5896 4494 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 4488 5868 5365 5896
rect 4488 5856 4494 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 5353 5859 5411 5865
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 5592 5868 8953 5896
rect 5592 5856 5598 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 10778 5896 10784 5908
rect 10739 5868 10784 5896
rect 8941 5859 8999 5865
rect 10778 5856 10784 5868
rect 10836 5856 10842 5908
rect 12802 5896 12808 5908
rect 12763 5868 12808 5896
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 3050 5828 3056 5840
rect 2056 5800 2774 5828
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 1854 5692 1860 5704
rect 1627 5664 1860 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 1854 5652 1860 5664
rect 1912 5652 1918 5704
rect 2056 5701 2084 5800
rect 2746 5704 2774 5800
rect 2884 5800 3056 5828
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2746 5664 2780 5704
rect 2225 5655 2283 5661
rect 2240 5624 2268 5655
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 2884 5701 2912 5800
rect 3050 5788 3056 5800
rect 3108 5788 3114 5840
rect 3234 5788 3240 5840
rect 3292 5788 3298 5840
rect 3252 5760 3280 5788
rect 2976 5732 3280 5760
rect 2976 5701 3004 5732
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5661 3019 5695
rect 2961 5655 3019 5661
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 4448 5692 4476 5856
rect 4801 5831 4859 5837
rect 4801 5797 4813 5831
rect 4847 5828 4859 5831
rect 5442 5828 5448 5840
rect 4847 5800 5448 5828
rect 4847 5797 4859 5800
rect 4801 5791 4859 5797
rect 5442 5788 5448 5800
rect 5500 5788 5506 5840
rect 5552 5760 5580 5856
rect 7006 5788 7012 5840
rect 7064 5828 7070 5840
rect 7064 5800 7144 5828
rect 7064 5788 7070 5800
rect 4908 5732 5580 5760
rect 7116 5760 7144 5800
rect 7650 5788 7656 5840
rect 7708 5828 7714 5840
rect 8113 5831 8171 5837
rect 7708 5800 8064 5828
rect 7708 5788 7714 5800
rect 7285 5763 7343 5769
rect 7285 5760 7297 5763
rect 7116 5732 7297 5760
rect 3283 5664 4476 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 4706 5701 4712 5704
rect 4677 5695 4712 5701
rect 4580 5664 4625 5692
rect 4580 5652 4586 5664
rect 4677 5661 4689 5695
rect 4677 5655 4712 5661
rect 4706 5652 4712 5655
rect 4764 5652 4770 5704
rect 4908 5701 4936 5732
rect 7285 5729 7297 5732
rect 7331 5729 7343 5763
rect 7926 5760 7932 5772
rect 7887 5732 7932 5760
rect 7285 5723 7343 5729
rect 7926 5720 7932 5732
rect 7984 5720 7990 5772
rect 8036 5769 8064 5800
rect 8113 5797 8125 5831
rect 8159 5828 8171 5831
rect 8202 5828 8208 5840
rect 8159 5800 8208 5828
rect 8159 5797 8171 5800
rect 8113 5791 8171 5797
rect 8202 5788 8208 5800
rect 8260 5788 8266 5840
rect 11241 5831 11299 5837
rect 11241 5828 11253 5831
rect 8312 5800 11253 5828
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5729 8079 5763
rect 8312 5760 8340 5800
rect 11241 5797 11253 5800
rect 11287 5797 11299 5831
rect 13354 5828 13360 5840
rect 13315 5800 13360 5828
rect 11241 5791 11299 5797
rect 13354 5788 13360 5800
rect 13412 5788 13418 5840
rect 14734 5788 14740 5840
rect 14792 5828 14798 5840
rect 14792 5800 15240 5828
rect 14792 5788 14798 5800
rect 9585 5763 9643 5769
rect 9585 5760 9597 5763
rect 8021 5723 8079 5729
rect 8128 5732 8340 5760
rect 9140 5732 9597 5760
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 5074 5652 5080 5704
rect 5132 5692 5138 5704
rect 5537 5695 5595 5701
rect 5537 5692 5549 5695
rect 5132 5664 5549 5692
rect 5132 5652 5138 5664
rect 5537 5661 5549 5664
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 5813 5695 5871 5701
rect 5813 5661 5825 5695
rect 5859 5692 5871 5695
rect 5902 5692 5908 5704
rect 5859 5664 5908 5692
rect 5859 5661 5871 5664
rect 5813 5655 5871 5661
rect 5902 5652 5908 5664
rect 5960 5692 5966 5704
rect 6641 5695 6699 5701
rect 6641 5692 6653 5695
rect 5960 5664 6653 5692
rect 5960 5652 5966 5664
rect 6641 5661 6653 5664
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 6730 5652 6736 5704
rect 6788 5691 6794 5704
rect 6825 5695 6883 5701
rect 6825 5691 6837 5695
rect 6788 5663 6837 5691
rect 6788 5652 6794 5663
rect 6825 5661 6837 5663
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 6917 5695 6975 5701
rect 6917 5661 6929 5695
rect 6963 5691 6975 5695
rect 7558 5692 7564 5704
rect 7116 5691 7564 5692
rect 6963 5664 7564 5691
rect 6963 5663 7144 5664
rect 6963 5661 6975 5663
rect 6917 5655 6975 5661
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5692 7803 5695
rect 8128 5692 8156 5732
rect 7791 5664 8156 5692
rect 8205 5695 8263 5701
rect 7791 5661 7803 5664
rect 7745 5655 7803 5661
rect 8205 5661 8217 5695
rect 8251 5692 8263 5695
rect 8294 5692 8300 5704
rect 8251 5664 8300 5692
rect 8251 5661 8263 5664
rect 8205 5655 8263 5661
rect 4062 5624 4068 5636
rect 2240 5596 4068 5624
rect 4062 5584 4068 5596
rect 4120 5584 4126 5636
rect 6454 5584 6460 5636
rect 6512 5624 6518 5636
rect 7009 5627 7067 5633
rect 7009 5624 7021 5627
rect 6512 5596 7021 5624
rect 6512 5584 6518 5596
rect 7009 5593 7021 5596
rect 7055 5593 7067 5627
rect 7009 5587 7067 5593
rect 7147 5627 7205 5633
rect 7147 5593 7159 5627
rect 7193 5624 7205 5627
rect 7466 5624 7472 5636
rect 7193 5596 7472 5624
rect 7193 5593 7205 5596
rect 7147 5587 7205 5593
rect 7466 5584 7472 5596
rect 7524 5584 7530 5636
rect 1394 5516 1400 5568
rect 1452 5556 1458 5568
rect 1489 5559 1547 5565
rect 1489 5556 1501 5559
rect 1452 5528 1501 5556
rect 1452 5516 1458 5528
rect 1489 5525 1501 5528
rect 1535 5525 1547 5559
rect 2130 5556 2136 5568
rect 2091 5528 2136 5556
rect 1489 5519 1547 5525
rect 2130 5516 2136 5528
rect 2188 5516 2194 5568
rect 2685 5559 2743 5565
rect 2685 5525 2697 5559
rect 2731 5556 2743 5559
rect 3418 5556 3424 5568
rect 2731 5528 3424 5556
rect 2731 5525 2743 5528
rect 2685 5519 2743 5525
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 5718 5556 5724 5568
rect 5679 5528 5724 5556
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 7760 5556 7788 5655
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 9140 5701 9168 5732
rect 9585 5729 9597 5732
rect 9631 5729 9643 5763
rect 9585 5723 9643 5729
rect 10229 5763 10287 5769
rect 10229 5729 10241 5763
rect 10275 5760 10287 5763
rect 11609 5763 11667 5769
rect 11609 5760 11621 5763
rect 10275 5732 11621 5760
rect 10275 5729 10287 5732
rect 10229 5723 10287 5729
rect 11609 5729 11621 5732
rect 11655 5760 11667 5763
rect 14826 5760 14832 5772
rect 11655 5732 12434 5760
rect 11655 5729 11667 5732
rect 11609 5723 11667 5729
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 8444 5664 9137 5692
rect 8444 5652 8450 5664
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 8478 5584 8484 5636
rect 8536 5624 8542 5636
rect 9232 5624 9260 5655
rect 9493 5627 9551 5633
rect 9493 5624 9505 5627
rect 8536 5596 9505 5624
rect 8536 5584 8542 5596
rect 9493 5593 9505 5596
rect 9539 5593 9551 5627
rect 9600 5624 9628 5723
rect 9858 5652 9864 5704
rect 9916 5692 9922 5704
rect 10505 5695 10563 5701
rect 9916 5691 10456 5692
rect 10505 5691 10517 5695
rect 9916 5664 10517 5691
rect 9916 5652 9922 5664
rect 10428 5663 10517 5664
rect 10505 5661 10517 5663
rect 10551 5661 10563 5695
rect 11425 5695 11483 5701
rect 11425 5692 11437 5695
rect 10505 5655 10563 5661
rect 10612 5664 11437 5692
rect 10612 5624 10640 5664
rect 11425 5661 11437 5664
rect 11471 5661 11483 5695
rect 11425 5655 11483 5661
rect 11514 5652 11520 5704
rect 11572 5692 11578 5704
rect 11701 5695 11759 5701
rect 11572 5664 11617 5692
rect 11572 5652 11578 5664
rect 11701 5661 11713 5695
rect 11747 5661 11759 5695
rect 12406 5692 12434 5732
rect 13924 5732 14832 5760
rect 13446 5692 13452 5704
rect 12406 5664 13452 5692
rect 11701 5655 11759 5661
rect 9600 5596 10640 5624
rect 9493 5587 9551 5593
rect 10962 5584 10968 5636
rect 11020 5624 11026 5636
rect 11716 5624 11744 5655
rect 13446 5652 13452 5664
rect 13504 5692 13510 5704
rect 13722 5692 13728 5704
rect 13504 5664 13728 5692
rect 13504 5652 13510 5664
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 11020 5596 11744 5624
rect 11020 5584 11026 5596
rect 12434 5584 12440 5636
rect 12492 5624 12498 5636
rect 13081 5627 13139 5633
rect 13081 5624 13093 5627
rect 12492 5596 13093 5624
rect 12492 5584 12498 5596
rect 13081 5593 13093 5596
rect 13127 5624 13139 5627
rect 13538 5624 13544 5636
rect 13127 5596 13544 5624
rect 13127 5593 13139 5596
rect 13081 5587 13139 5593
rect 13538 5584 13544 5596
rect 13596 5584 13602 5636
rect 6604 5528 7788 5556
rect 6604 5516 6610 5528
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 8389 5559 8447 5565
rect 8389 5556 8401 5559
rect 8260 5528 8401 5556
rect 8260 5516 8266 5528
rect 8389 5525 8401 5528
rect 8435 5525 8447 5559
rect 10410 5556 10416 5568
rect 10371 5528 10416 5556
rect 8389 5519 8447 5525
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 10502 5516 10508 5568
rect 10560 5556 10566 5568
rect 10597 5559 10655 5565
rect 10597 5556 10609 5559
rect 10560 5528 10609 5556
rect 10560 5516 10566 5528
rect 10597 5525 10609 5528
rect 10643 5525 10655 5559
rect 10597 5519 10655 5525
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 12158 5556 12164 5568
rect 10744 5528 12164 5556
rect 10744 5516 10750 5528
rect 12158 5516 12164 5528
rect 12216 5516 12222 5568
rect 12342 5516 12348 5568
rect 12400 5556 12406 5568
rect 12986 5556 12992 5568
rect 12400 5528 12992 5556
rect 12400 5516 12406 5528
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 13173 5559 13231 5565
rect 13173 5525 13185 5559
rect 13219 5556 13231 5559
rect 13924 5556 13952 5732
rect 14826 5720 14832 5732
rect 14884 5720 14890 5772
rect 15010 5760 15016 5772
rect 14971 5732 15016 5760
rect 15010 5720 15016 5732
rect 15068 5720 15074 5772
rect 15212 5760 15240 5800
rect 15212 5732 15332 5760
rect 14366 5652 14372 5704
rect 14424 5692 14430 5704
rect 14461 5695 14519 5701
rect 14461 5692 14473 5695
rect 14424 5664 14473 5692
rect 14424 5652 14430 5664
rect 14461 5661 14473 5664
rect 14507 5661 14519 5695
rect 14461 5655 14519 5661
rect 14550 5652 14556 5704
rect 14608 5692 14614 5704
rect 14921 5695 14979 5701
rect 14921 5692 14933 5695
rect 14608 5664 14933 5692
rect 14608 5652 14614 5664
rect 14921 5661 14933 5664
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 15102 5652 15108 5704
rect 15160 5692 15166 5704
rect 15304 5701 15332 5732
rect 15197 5695 15255 5701
rect 15197 5692 15209 5695
rect 15160 5664 15209 5692
rect 15160 5652 15166 5664
rect 15197 5661 15209 5664
rect 15243 5661 15255 5695
rect 15197 5655 15255 5661
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 14277 5627 14335 5633
rect 14277 5593 14289 5627
rect 14323 5624 14335 5627
rect 14642 5624 14648 5636
rect 14323 5596 14648 5624
rect 14323 5593 14335 5596
rect 14277 5587 14335 5593
rect 14642 5584 14648 5596
rect 14700 5584 14706 5636
rect 15212 5624 15240 5655
rect 15378 5624 15384 5636
rect 15212 5596 15384 5624
rect 15378 5584 15384 5596
rect 15436 5584 15442 5636
rect 14090 5556 14096 5568
rect 13219 5528 13952 5556
rect 14051 5528 14096 5556
rect 13219 5525 13231 5528
rect 13173 5519 13231 5525
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 15473 5559 15531 5565
rect 15473 5556 15485 5559
rect 15252 5528 15485 5556
rect 15252 5516 15258 5528
rect 15473 5525 15485 5528
rect 15519 5525 15531 5559
rect 15473 5519 15531 5525
rect 1104 5466 16468 5488
rect 1104 5414 6103 5466
rect 6155 5414 6167 5466
rect 6219 5414 6231 5466
rect 6283 5414 6295 5466
rect 6347 5414 11224 5466
rect 11276 5414 11288 5466
rect 11340 5414 11352 5466
rect 11404 5414 11416 5466
rect 11468 5414 16468 5466
rect 1104 5392 16468 5414
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 3326 5352 3332 5364
rect 2832 5324 3332 5352
rect 2832 5312 2838 5324
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 3881 5355 3939 5361
rect 3881 5321 3893 5355
rect 3927 5321 3939 5355
rect 3881 5315 3939 5321
rect 3237 5287 3295 5293
rect 3237 5253 3249 5287
rect 3283 5284 3295 5287
rect 3896 5284 3924 5315
rect 6730 5312 6736 5364
rect 6788 5352 6794 5364
rect 7558 5352 7564 5364
rect 6788 5324 7564 5352
rect 6788 5312 6794 5324
rect 7558 5312 7564 5324
rect 7616 5352 7622 5364
rect 8202 5352 8208 5364
rect 7616 5324 8208 5352
rect 7616 5312 7622 5324
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 10410 5352 10416 5364
rect 10371 5324 10416 5352
rect 10410 5312 10416 5324
rect 10468 5312 10474 5364
rect 10502 5312 10508 5364
rect 10560 5352 10566 5364
rect 12434 5352 12440 5364
rect 10560 5324 10605 5352
rect 10704 5324 12440 5352
rect 10560 5312 10566 5324
rect 3970 5284 3976 5296
rect 3283 5256 3976 5284
rect 3283 5253 3295 5256
rect 3237 5247 3295 5253
rect 3970 5244 3976 5256
rect 4028 5244 4034 5296
rect 4525 5287 4583 5293
rect 4525 5284 4537 5287
rect 4080 5256 4537 5284
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 1762 5216 1768 5228
rect 1719 5188 1768 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 1762 5176 1768 5188
rect 1820 5176 1826 5228
rect 2314 5216 2320 5228
rect 2275 5188 2320 5216
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 3418 5216 3424 5228
rect 3379 5188 3424 5216
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 4080 5225 4108 5256
rect 4525 5253 4537 5256
rect 4571 5253 4583 5287
rect 4525 5247 4583 5253
rect 5074 5244 5080 5296
rect 5132 5284 5138 5296
rect 5353 5287 5411 5293
rect 5353 5284 5365 5287
rect 5132 5256 5365 5284
rect 5132 5244 5138 5256
rect 5353 5253 5365 5256
rect 5399 5253 5411 5287
rect 5353 5247 5411 5253
rect 6932 5256 8984 5284
rect 6932 5228 6960 5256
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 5166 5216 5172 5228
rect 4203 5188 4476 5216
rect 5127 5188 5172 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 4080 5080 4108 5179
rect 4448 5157 4476 5188
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5216 5319 5219
rect 5534 5216 5540 5228
rect 5307 5188 5396 5216
rect 5495 5188 5540 5216
rect 5307 5185 5319 5188
rect 5261 5179 5319 5185
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 4479 5120 5120 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 4982 5080 4988 5092
rect 4080 5052 4988 5080
rect 4982 5040 4988 5052
rect 5040 5040 5046 5092
rect 5092 5024 5120 5120
rect 5368 5092 5396 5188
rect 5534 5176 5540 5188
rect 5592 5176 5598 5228
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 6914 5216 6920 5228
rect 5684 5188 6920 5216
rect 5684 5176 5690 5188
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 7064 5188 7205 5216
rect 7064 5176 7070 5188
rect 7193 5185 7205 5188
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 7466 5216 7472 5228
rect 7423 5188 7472 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 7834 5216 7840 5228
rect 7795 5188 7840 5216
rect 7834 5176 7840 5188
rect 7892 5176 7898 5228
rect 8956 5225 8984 5256
rect 9858 5244 9864 5296
rect 9916 5284 9922 5296
rect 10229 5287 10287 5293
rect 10229 5284 10241 5287
rect 9916 5256 10241 5284
rect 9916 5244 9922 5256
rect 10229 5253 10241 5256
rect 10275 5284 10287 5287
rect 10704 5284 10732 5324
rect 12434 5312 12440 5324
rect 12492 5312 12498 5364
rect 12894 5352 12900 5364
rect 12855 5324 12900 5352
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 13538 5312 13544 5364
rect 13596 5352 13602 5364
rect 14185 5355 14243 5361
rect 14185 5352 14197 5355
rect 13596 5324 14197 5352
rect 13596 5312 13602 5324
rect 14185 5321 14197 5324
rect 14231 5321 14243 5355
rect 14185 5315 14243 5321
rect 14461 5355 14519 5361
rect 14461 5321 14473 5355
rect 14507 5352 14519 5355
rect 14918 5352 14924 5364
rect 14507 5324 14924 5352
rect 14507 5321 14519 5324
rect 14461 5315 14519 5321
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 12805 5287 12863 5293
rect 12805 5284 12817 5287
rect 10275 5256 10732 5284
rect 11808 5256 12817 5284
rect 10275 5253 10287 5256
rect 10229 5247 10287 5253
rect 11808 5228 11836 5256
rect 12805 5253 12817 5256
rect 12851 5253 12863 5287
rect 12805 5247 12863 5253
rect 12912 5256 13768 5284
rect 8941 5219 8999 5225
rect 8941 5185 8953 5219
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 11790 5216 11796 5228
rect 10652 5188 10697 5216
rect 11703 5188 11796 5216
rect 10652 5176 10658 5188
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5216 11943 5219
rect 11974 5216 11980 5228
rect 11931 5188 11980 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5216 12219 5219
rect 12434 5216 12440 5228
rect 12207 5188 12440 5216
rect 12207 5185 12219 5188
rect 12161 5179 12219 5185
rect 12434 5176 12440 5188
rect 12492 5176 12498 5228
rect 12912 5216 12940 5256
rect 12728 5188 12940 5216
rect 13081 5219 13139 5225
rect 6638 5108 6644 5160
rect 6696 5148 6702 5160
rect 7101 5151 7159 5157
rect 7101 5148 7113 5151
rect 6696 5120 7113 5148
rect 6696 5108 6702 5120
rect 7101 5117 7113 5120
rect 7147 5148 7159 5151
rect 7650 5148 7656 5160
rect 7147 5120 7656 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 8665 5151 8723 5157
rect 8665 5148 8677 5151
rect 8352 5120 8677 5148
rect 8352 5108 8358 5120
rect 8665 5117 8677 5120
rect 8711 5148 8723 5151
rect 10686 5148 10692 5160
rect 8711 5120 10692 5148
rect 8711 5117 8723 5120
rect 8665 5111 8723 5117
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 11606 5108 11612 5160
rect 11664 5108 11670 5160
rect 11698 5108 11704 5160
rect 11756 5148 11762 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11756 5120 12081 5148
rect 11756 5108 11762 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 5350 5040 5356 5092
rect 5408 5040 5414 5092
rect 6822 5040 6828 5092
rect 6880 5080 6886 5092
rect 7009 5083 7067 5089
rect 7009 5080 7021 5083
rect 6880 5052 7021 5080
rect 6880 5040 6886 5052
rect 7009 5049 7021 5052
rect 7055 5080 7067 5083
rect 8202 5080 8208 5092
rect 7055 5052 8208 5080
rect 7055 5049 7067 5052
rect 7009 5043 7067 5049
rect 8202 5040 8208 5052
rect 8260 5040 8266 5092
rect 10962 5080 10968 5092
rect 10796 5052 10968 5080
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 1670 4972 1676 5024
rect 1728 5012 1734 5024
rect 2225 5015 2283 5021
rect 2225 5012 2237 5015
rect 1728 4984 2237 5012
rect 1728 4972 1734 4984
rect 2225 4981 2237 4984
rect 2271 4981 2283 5015
rect 2225 4975 2283 4981
rect 2866 4972 2872 5024
rect 2924 5012 2930 5024
rect 3053 5015 3111 5021
rect 3053 5012 3065 5015
rect 2924 4984 3065 5012
rect 2924 4972 2930 4984
rect 3053 4981 3065 4984
rect 3099 4981 3111 5015
rect 3053 4975 3111 4981
rect 5074 4972 5080 5024
rect 5132 5012 5138 5024
rect 6733 5015 6791 5021
rect 6733 5012 6745 5015
rect 5132 4984 6745 5012
rect 5132 4972 5138 4984
rect 6733 4981 6745 4984
rect 6779 4981 6791 5015
rect 8018 5012 8024 5024
rect 7979 4984 8024 5012
rect 6733 4975 6791 4981
rect 8018 4972 8024 4984
rect 8076 4972 8082 5024
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 10796 5021 10824 5052
rect 10962 5040 10968 5052
rect 11020 5040 11026 5092
rect 11624 5080 11652 5108
rect 12250 5080 12256 5092
rect 11624 5052 12256 5080
rect 12250 5040 12256 5052
rect 12308 5080 12314 5092
rect 12308 5052 12434 5080
rect 12308 5040 12314 5052
rect 10781 5015 10839 5021
rect 10781 5012 10793 5015
rect 8352 4984 10793 5012
rect 8352 4972 8358 4984
rect 10781 4981 10793 4984
rect 10827 4981 10839 5015
rect 10781 4975 10839 4981
rect 10870 4972 10876 5024
rect 10928 5012 10934 5024
rect 11609 5015 11667 5021
rect 11609 5012 11621 5015
rect 10928 4984 11621 5012
rect 10928 4972 10934 4984
rect 11609 4981 11621 4984
rect 11655 4981 11667 5015
rect 12406 5012 12434 5052
rect 12728 5012 12756 5188
rect 13081 5185 13093 5219
rect 13127 5185 13139 5219
rect 13081 5179 13139 5185
rect 13173 5219 13231 5225
rect 13173 5185 13185 5219
rect 13219 5185 13231 5219
rect 13173 5179 13231 5185
rect 13449 5219 13507 5225
rect 13449 5185 13461 5219
rect 13495 5216 13507 5219
rect 13495 5188 13676 5216
rect 13495 5185 13507 5188
rect 13449 5179 13507 5185
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5148 12863 5151
rect 12894 5148 12900 5160
rect 12851 5120 12900 5148
rect 12851 5117 12863 5120
rect 12805 5111 12863 5117
rect 12894 5108 12900 5120
rect 12952 5148 12958 5160
rect 13096 5148 13124 5179
rect 12952 5120 13124 5148
rect 12952 5108 12958 5120
rect 12406 4984 12756 5012
rect 13188 5012 13216 5179
rect 13354 5108 13360 5160
rect 13412 5148 13418 5160
rect 13412 5120 13457 5148
rect 13412 5108 13418 5120
rect 13648 5080 13676 5188
rect 13740 5148 13768 5256
rect 13906 5244 13912 5296
rect 13964 5284 13970 5296
rect 13964 5256 14009 5284
rect 13964 5244 13970 5256
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 13872 5188 14105 5216
rect 13872 5176 13878 5188
rect 14093 5185 14105 5188
rect 14139 5185 14151 5219
rect 14093 5179 14151 5185
rect 14277 5219 14335 5225
rect 14277 5185 14289 5219
rect 14323 5216 14335 5219
rect 15102 5216 15108 5228
rect 14323 5188 15108 5216
rect 14323 5185 14335 5188
rect 14277 5179 14335 5185
rect 14292 5148 14320 5179
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 13740 5120 14320 5148
rect 14550 5108 14556 5160
rect 14608 5148 14614 5160
rect 14921 5151 14979 5157
rect 14921 5148 14933 5151
rect 14608 5120 14933 5148
rect 14608 5108 14614 5120
rect 14921 5117 14933 5120
rect 14967 5117 14979 5151
rect 14921 5111 14979 5117
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5148 15255 5151
rect 16669 5151 16727 5157
rect 16669 5148 16681 5151
rect 15243 5120 16681 5148
rect 15243 5117 15255 5120
rect 15197 5111 15255 5117
rect 16669 5117 16681 5120
rect 16715 5117 16727 5151
rect 16669 5111 16727 5117
rect 15212 5080 15240 5111
rect 13648 5052 15240 5080
rect 14182 5012 14188 5024
rect 13188 4984 14188 5012
rect 11609 4975 11667 4981
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 1104 4922 16468 4944
rect 1104 4870 3542 4922
rect 3594 4870 3606 4922
rect 3658 4870 3670 4922
rect 3722 4870 3734 4922
rect 3786 4870 8664 4922
rect 8716 4870 8728 4922
rect 8780 4870 8792 4922
rect 8844 4870 8856 4922
rect 8908 4870 13785 4922
rect 13837 4870 13849 4922
rect 13901 4870 13913 4922
rect 13965 4870 13977 4922
rect 14029 4870 16468 4922
rect 1104 4848 16468 4870
rect 1578 4768 1584 4820
rect 1636 4808 1642 4820
rect 1765 4811 1823 4817
rect 1765 4808 1777 4811
rect 1636 4780 1777 4808
rect 1636 4768 1642 4780
rect 1765 4777 1777 4780
rect 1811 4777 1823 4811
rect 1765 4771 1823 4777
rect 3145 4811 3203 4817
rect 3145 4777 3157 4811
rect 3191 4808 3203 4811
rect 5166 4808 5172 4820
rect 3191 4780 5172 4808
rect 3191 4777 3203 4780
rect 3145 4771 3203 4777
rect 5166 4768 5172 4780
rect 5224 4808 5230 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 5224 4780 5273 4808
rect 5224 4768 5230 4780
rect 5261 4777 5273 4780
rect 5307 4777 5319 4811
rect 5261 4771 5319 4777
rect 7285 4811 7343 4817
rect 7285 4777 7297 4811
rect 7331 4808 7343 4811
rect 7834 4808 7840 4820
rect 7331 4780 7840 4808
rect 7331 4777 7343 4780
rect 7285 4771 7343 4777
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 8386 4808 8392 4820
rect 8347 4780 8392 4808
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 10134 4768 10140 4820
rect 10192 4808 10198 4820
rect 10413 4811 10471 4817
rect 10413 4808 10425 4811
rect 10192 4780 10425 4808
rect 10192 4768 10198 4780
rect 10413 4777 10425 4780
rect 10459 4777 10471 4811
rect 11698 4808 11704 4820
rect 11659 4780 11704 4808
rect 10413 4771 10471 4777
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 13170 4808 13176 4820
rect 13131 4780 13176 4808
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 13354 4808 13360 4820
rect 13315 4780 13360 4808
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 14093 4811 14151 4817
rect 14093 4777 14105 4811
rect 14139 4808 14151 4811
rect 14182 4808 14188 4820
rect 14139 4780 14188 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 4798 4740 4804 4752
rect 3252 4712 4804 4740
rect 1670 4604 1676 4616
rect 1631 4576 1676 4604
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 1762 4564 1768 4616
rect 1820 4604 1826 4616
rect 1946 4604 1952 4616
rect 1820 4576 1952 4604
rect 1820 4564 1826 4576
rect 1946 4564 1952 4576
rect 2004 4564 2010 4616
rect 3252 4613 3280 4712
rect 4798 4700 4804 4712
rect 4856 4740 4862 4752
rect 5442 4740 5448 4752
rect 4856 4712 5448 4740
rect 4856 4700 4862 4712
rect 5442 4700 5448 4712
rect 5500 4700 5506 4752
rect 3418 4632 3424 4684
rect 3476 4672 3482 4684
rect 3789 4675 3847 4681
rect 3789 4672 3801 4675
rect 3476 4644 3801 4672
rect 3476 4632 3482 4644
rect 3789 4641 3801 4644
rect 3835 4641 3847 4675
rect 11241 4675 11299 4681
rect 11241 4672 11253 4675
rect 3789 4635 3847 4641
rect 8220 4644 11253 4672
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4573 2099 4607
rect 2041 4567 2099 4573
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4573 3295 4607
rect 3970 4604 3976 4616
rect 3931 4576 3976 4604
rect 3237 4567 3295 4573
rect 2056 4536 2084 4567
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 4338 4604 4344 4616
rect 4299 4576 4344 4604
rect 4338 4564 4344 4576
rect 4396 4564 4402 4616
rect 4982 4604 4988 4616
rect 4943 4576 4988 4604
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 5074 4564 5080 4616
rect 5132 4604 5138 4616
rect 5350 4604 5356 4616
rect 5132 4576 5177 4604
rect 5311 4576 5356 4604
rect 5132 4564 5138 4576
rect 5350 4564 5356 4576
rect 5408 4604 5414 4616
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 5408 4576 5825 4604
rect 5408 4564 5414 4576
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 5902 4564 5908 4616
rect 5960 4604 5966 4616
rect 6181 4607 6239 4613
rect 6181 4604 6193 4607
rect 5960 4576 6193 4604
rect 5960 4564 5966 4576
rect 6181 4573 6193 4576
rect 6227 4573 6239 4607
rect 7190 4604 7196 4616
rect 7151 4576 7196 4604
rect 6181 4567 6239 4573
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 8220 4613 8248 4644
rect 11241 4641 11253 4644
rect 11287 4641 11299 4675
rect 11716 4672 11744 4768
rect 13262 4700 13268 4752
rect 13320 4740 13326 4752
rect 13538 4740 13544 4752
rect 13320 4712 13544 4740
rect 13320 4700 13326 4712
rect 13538 4700 13544 4712
rect 13596 4700 13602 4752
rect 13449 4675 13507 4681
rect 11241 4635 11299 4641
rect 11440 4644 11652 4672
rect 11716 4644 12388 4672
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 8389 4607 8447 4613
rect 8389 4604 8401 4607
rect 8352 4576 8401 4604
rect 8352 4564 8358 4576
rect 8389 4573 8401 4576
rect 8435 4573 8447 4607
rect 8938 4604 8944 4616
rect 8899 4576 8944 4604
rect 8389 4567 8447 4573
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 9214 4604 9220 4616
rect 9175 4576 9220 4604
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4604 10655 4607
rect 10870 4604 10876 4616
rect 10643 4576 10876 4604
rect 10643 4573 10655 4576
rect 10597 4567 10655 4573
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 11440 4613 11468 4644
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4573 11483 4607
rect 11425 4567 11483 4573
rect 11517 4607 11575 4613
rect 11517 4573 11529 4607
rect 11563 4573 11575 4607
rect 11517 4567 11575 4573
rect 2314 4536 2320 4548
rect 2056 4508 2320 4536
rect 2314 4496 2320 4508
rect 2372 4536 2378 4548
rect 2372 4508 4016 4536
rect 2372 4496 2378 4508
rect 2225 4471 2283 4477
rect 2225 4437 2237 4471
rect 2271 4468 2283 4471
rect 2958 4468 2964 4480
rect 2271 4440 2964 4468
rect 2271 4437 2283 4440
rect 2225 4431 2283 4437
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 3988 4477 4016 4508
rect 4062 4496 4068 4548
rect 4120 4536 4126 4548
rect 4801 4539 4859 4545
rect 4801 4536 4813 4539
rect 4120 4508 4813 4536
rect 4120 4496 4126 4508
rect 4801 4505 4813 4508
rect 4847 4505 4859 4539
rect 4801 4499 4859 4505
rect 5718 4496 5724 4548
rect 5776 4536 5782 4548
rect 5997 4539 6055 4545
rect 5997 4536 6009 4539
rect 5776 4508 6009 4536
rect 5776 4496 5782 4508
rect 5997 4505 6009 4508
rect 6043 4536 6055 4539
rect 9306 4536 9312 4548
rect 6043 4508 9312 4536
rect 6043 4505 6055 4508
rect 5997 4499 6055 4505
rect 9306 4496 9312 4508
rect 9364 4496 9370 4548
rect 10778 4536 10784 4548
rect 10739 4508 10784 4536
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 11054 4496 11060 4548
rect 11112 4536 11118 4548
rect 11532 4536 11560 4567
rect 11112 4508 11560 4536
rect 11624 4536 11652 4644
rect 11790 4604 11796 4616
rect 11751 4576 11796 4604
rect 11790 4564 11796 4576
rect 11848 4564 11854 4616
rect 12360 4613 12388 4644
rect 13449 4641 13461 4675
rect 13495 4672 13507 4675
rect 14108 4672 14136 4771
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 13495 4644 14136 4672
rect 14829 4675 14887 4681
rect 13495 4641 13507 4644
rect 13449 4635 13507 4641
rect 14829 4641 14841 4675
rect 14875 4672 14887 4675
rect 15010 4672 15016 4684
rect 14875 4644 15016 4672
rect 14875 4641 14887 4644
rect 14829 4635 14887 4641
rect 15010 4632 15016 4644
rect 15068 4632 15074 4684
rect 12345 4607 12403 4613
rect 12345 4573 12357 4607
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 13538 4564 13544 4616
rect 13596 4604 13602 4616
rect 14277 4607 14335 4613
rect 13596 4576 13641 4604
rect 13596 4564 13602 4576
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 14366 4604 14372 4616
rect 14323 4576 14372 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 14642 4564 14648 4616
rect 14700 4604 14706 4616
rect 15105 4607 15163 4613
rect 15105 4604 15117 4607
rect 14700 4576 15117 4604
rect 14700 4564 14706 4576
rect 15105 4573 15117 4576
rect 15151 4573 15163 4607
rect 15105 4567 15163 4573
rect 11974 4536 11980 4548
rect 11624 4508 11980 4536
rect 11112 4496 11118 4508
rect 11974 4496 11980 4508
rect 12032 4496 12038 4548
rect 12529 4539 12587 4545
rect 12529 4505 12541 4539
rect 12575 4536 12587 4539
rect 12710 4536 12716 4548
rect 12575 4508 12716 4536
rect 12575 4505 12587 4508
rect 12529 4499 12587 4505
rect 12710 4496 12716 4508
rect 12768 4496 12774 4548
rect 12894 4496 12900 4548
rect 12952 4536 12958 4548
rect 14734 4536 14740 4548
rect 12952 4508 14740 4536
rect 12952 4496 12958 4508
rect 14734 4496 14740 4508
rect 14792 4496 14798 4548
rect 3973 4471 4031 4477
rect 3973 4437 3985 4471
rect 4019 4437 4031 4471
rect 3973 4431 4031 4437
rect 5166 4428 5172 4480
rect 5224 4468 5230 4480
rect 8110 4468 8116 4480
rect 5224 4440 8116 4468
rect 5224 4428 5230 4440
rect 8110 4428 8116 4440
rect 8168 4468 8174 4480
rect 8938 4468 8944 4480
rect 8168 4440 8944 4468
rect 8168 4428 8174 4440
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 15010 4468 15016 4480
rect 12492 4440 15016 4468
rect 12492 4428 12498 4440
rect 15010 4428 15016 4440
rect 15068 4428 15074 4480
rect 1104 4378 16468 4400
rect 1104 4326 6103 4378
rect 6155 4326 6167 4378
rect 6219 4326 6231 4378
rect 6283 4326 6295 4378
rect 6347 4326 11224 4378
rect 11276 4326 11288 4378
rect 11340 4326 11352 4378
rect 11404 4326 11416 4378
rect 11468 4326 16468 4378
rect 1104 4304 16468 4326
rect 4522 4264 4528 4276
rect 4080 4236 4528 4264
rect 1670 4128 1676 4140
rect 1631 4100 1676 4128
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 2866 4128 2872 4140
rect 2746 4100 2872 4128
rect 1578 4020 1584 4072
rect 1636 4060 1642 4072
rect 1765 4063 1823 4069
rect 1765 4060 1777 4063
rect 1636 4032 1777 4060
rect 1636 4020 1642 4032
rect 1765 4029 1777 4032
rect 1811 4029 1823 4063
rect 1765 4023 1823 4029
rect 1949 4063 2007 4069
rect 1949 4029 1961 4063
rect 1995 4060 2007 4063
rect 2746 4060 2774 4100
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 4080 4128 4108 4236
rect 4522 4224 4528 4236
rect 4580 4224 4586 4276
rect 4890 4264 4896 4276
rect 4851 4236 4896 4264
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 8018 4264 8024 4276
rect 5368 4236 8024 4264
rect 5368 4196 5396 4236
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 8849 4267 8907 4273
rect 8849 4233 8861 4267
rect 8895 4233 8907 4267
rect 8849 4227 8907 4233
rect 4908 4168 5396 4196
rect 5445 4199 5503 4205
rect 3743 4100 4108 4128
rect 4157 4131 4215 4137
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 4157 4097 4169 4131
rect 4203 4126 4215 4131
rect 4908 4128 4936 4168
rect 5445 4165 5457 4199
rect 5491 4165 5503 4199
rect 7834 4196 7840 4208
rect 5445 4159 5503 4165
rect 6932 4168 7840 4196
rect 4264 4126 4936 4128
rect 4203 4100 4936 4126
rect 4985 4131 5043 4137
rect 4203 4098 4292 4100
rect 4203 4097 4215 4098
rect 4157 4091 4215 4097
rect 4985 4097 4997 4131
rect 5031 4128 5043 4131
rect 5350 4128 5356 4140
rect 5031 4100 5356 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5460 4072 5488 4159
rect 6932 4140 6960 4168
rect 7834 4156 7840 4168
rect 7892 4156 7898 4208
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 6730 4128 6736 4140
rect 5767 4100 6736 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 1995 4032 2774 4060
rect 2961 4063 3019 4069
rect 1995 4029 2007 4032
rect 1949 4023 2007 4029
rect 2961 4029 2973 4063
rect 3007 4060 3019 4063
rect 4338 4060 4344 4072
rect 3007 4032 4344 4060
rect 3007 4029 3019 4032
rect 2961 4023 3019 4029
rect 4338 4020 4344 4032
rect 4396 4020 4402 4072
rect 5442 4060 5448 4072
rect 5355 4032 5448 4060
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5644 4060 5672 4091
rect 6730 4088 6736 4100
rect 6788 4088 6794 4140
rect 6914 4128 6920 4140
rect 6875 4100 6920 4128
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7098 4128 7104 4140
rect 7059 4100 7104 4128
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 7190 4088 7196 4140
rect 7248 4128 7254 4140
rect 7561 4131 7619 4137
rect 7561 4128 7573 4131
rect 7248 4100 7573 4128
rect 7248 4088 7254 4100
rect 7561 4097 7573 4100
rect 7607 4097 7619 4131
rect 8864 4128 8892 4227
rect 12434 4224 12440 4276
rect 12492 4264 12498 4276
rect 12529 4267 12587 4273
rect 12529 4264 12541 4267
rect 12492 4236 12541 4264
rect 12492 4224 12498 4236
rect 12529 4233 12541 4236
rect 12575 4233 12587 4267
rect 12529 4227 12587 4233
rect 15286 4224 15292 4276
rect 15344 4264 15350 4276
rect 15381 4267 15439 4273
rect 15381 4264 15393 4267
rect 15344 4236 15393 4264
rect 15344 4224 15350 4236
rect 15381 4233 15393 4236
rect 15427 4233 15439 4267
rect 15381 4227 15439 4233
rect 9214 4156 9220 4208
rect 9272 4196 9278 4208
rect 10321 4199 10379 4205
rect 10321 4196 10333 4199
rect 9272 4168 10333 4196
rect 9272 4156 9278 4168
rect 10321 4165 10333 4168
rect 10367 4165 10379 4199
rect 12710 4196 12716 4208
rect 10321 4159 10379 4165
rect 11900 4168 12716 4196
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 7561 4091 7619 4097
rect 7668 4100 8892 4128
rect 8956 4100 9137 4128
rect 6822 4060 6828 4072
rect 5644 4032 6828 4060
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 7668 4060 7696 4100
rect 6932 4032 7696 4060
rect 3605 3995 3663 4001
rect 3605 3961 3617 3995
rect 3651 3992 3663 3995
rect 5460 3992 5488 4020
rect 6932 4004 6960 4032
rect 7742 4020 7748 4072
rect 7800 4060 7806 4072
rect 8956 4071 8984 4100
rect 9125 4097 9137 4100
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9456 4100 10057 4128
rect 9456 4088 9462 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10778 4128 10784 4140
rect 10739 4100 10784 4128
rect 10045 4091 10103 4097
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 11900 4128 11928 4168
rect 12452 4140 12480 4168
rect 12710 4156 12716 4168
rect 12768 4156 12774 4208
rect 14366 4196 14372 4208
rect 14327 4168 14372 4196
rect 14366 4156 14372 4168
rect 14424 4156 14430 4208
rect 14550 4196 14556 4208
rect 14511 4168 14556 4196
rect 14550 4156 14556 4168
rect 14608 4156 14614 4208
rect 14918 4156 14924 4208
rect 14976 4196 14982 4208
rect 15013 4199 15071 4205
rect 15013 4196 15025 4199
rect 14976 4168 15025 4196
rect 14976 4156 14982 4168
rect 15013 4165 15025 4168
rect 15059 4165 15071 4199
rect 15194 4196 15200 4208
rect 15155 4168 15200 4196
rect 15013 4159 15071 4165
rect 15194 4156 15200 4168
rect 15252 4156 15258 4208
rect 11747 4100 11928 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 11974 4088 11980 4140
rect 12032 4128 12038 4140
rect 12032 4100 12077 4128
rect 12032 4088 12038 4100
rect 12434 4088 12440 4140
rect 12492 4088 12498 4140
rect 12526 4088 12532 4140
rect 12584 4128 12590 4140
rect 12621 4131 12679 4137
rect 12621 4128 12633 4131
rect 12584 4100 12633 4128
rect 12584 4088 12590 4100
rect 12621 4097 12633 4100
rect 12667 4097 12679 4131
rect 12621 4091 12679 4097
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 13173 4131 13231 4137
rect 13173 4128 13185 4131
rect 13044 4100 13185 4128
rect 13044 4088 13050 4100
rect 13173 4097 13185 4100
rect 13219 4097 13231 4131
rect 13173 4091 13231 4097
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 14274 4128 14280 4140
rect 13311 4100 14280 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 7800 4032 7849 4060
rect 7800 4020 7806 4032
rect 7837 4029 7849 4032
rect 7883 4060 7895 4063
rect 8864 4060 8984 4071
rect 7883 4043 8984 4060
rect 9033 4063 9091 4069
rect 7883 4032 8892 4043
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 9033 4029 9045 4063
rect 9079 4029 9091 4063
rect 9033 4023 9091 4029
rect 9218 4063 9276 4069
rect 9218 4029 9230 4063
rect 9264 4029 9276 4063
rect 9218 4023 9276 4029
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 9490 4060 9496 4072
rect 9355 4032 9496 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 3651 3964 5488 3992
rect 3651 3961 3663 3964
rect 3605 3955 3663 3961
rect 6086 3952 6092 4004
rect 6144 3992 6150 4004
rect 6914 3992 6920 4004
rect 6144 3964 6920 3992
rect 6144 3952 6150 3964
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 7101 3995 7159 4001
rect 7101 3961 7113 3995
rect 7147 3992 7159 3995
rect 8478 3992 8484 4004
rect 7147 3964 8484 3992
rect 7147 3961 7159 3964
rect 7101 3955 7159 3961
rect 8478 3952 8484 3964
rect 8536 3952 8542 4004
rect 1762 3884 1768 3936
rect 1820 3924 1826 3936
rect 1857 3927 1915 3933
rect 1857 3924 1869 3927
rect 1820 3896 1869 3924
rect 1820 3884 1826 3896
rect 1857 3893 1869 3896
rect 1903 3893 1915 3927
rect 1857 3887 1915 3893
rect 4341 3927 4399 3933
rect 4341 3893 4353 3927
rect 4387 3924 4399 3927
rect 4706 3924 4712 3936
rect 4387 3896 4712 3924
rect 4387 3893 4399 3896
rect 4341 3887 4399 3893
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 4798 3884 4804 3936
rect 4856 3924 4862 3936
rect 5445 3927 5503 3933
rect 5445 3924 5457 3927
rect 4856 3896 5457 3924
rect 4856 3884 4862 3896
rect 5445 3893 5457 3896
rect 5491 3893 5503 3927
rect 5445 3887 5503 3893
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 9048 3924 9076 4023
rect 9232 3992 9260 4023
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 11793 4063 11851 4069
rect 11793 4060 11805 4063
rect 10275 4032 11805 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 11793 4029 11805 4032
rect 11839 4060 11851 4063
rect 12710 4060 12716 4072
rect 11839 4032 12716 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 14826 4060 14832 4072
rect 12820 4032 14832 4060
rect 10778 3992 10784 4004
rect 9232 3964 10784 3992
rect 10778 3952 10784 3964
rect 10836 3992 10842 4004
rect 12820 3992 12848 4032
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 10836 3964 12848 3992
rect 10836 3952 10842 3964
rect 12894 3952 12900 4004
rect 12952 3992 12958 4004
rect 13446 3992 13452 4004
rect 12952 3964 13452 3992
rect 12952 3952 12958 3964
rect 13446 3952 13452 3964
rect 13504 3992 13510 4004
rect 14458 3992 14464 4004
rect 13504 3964 14464 3992
rect 13504 3952 13510 3964
rect 14458 3952 14464 3964
rect 14516 3952 14522 4004
rect 8076 3896 9076 3924
rect 8076 3884 8082 3896
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 9861 3927 9919 3933
rect 9861 3924 9873 3927
rect 9732 3896 9873 3924
rect 9732 3884 9738 3896
rect 9861 3893 9873 3896
rect 9907 3893 9919 3927
rect 10318 3924 10324 3936
rect 10279 3896 10324 3924
rect 9861 3887 9919 3893
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 10873 3927 10931 3933
rect 10873 3893 10885 3927
rect 10919 3924 10931 3927
rect 11054 3924 11060 3936
rect 10919 3896 11060 3924
rect 10919 3893 10931 3896
rect 10873 3887 10931 3893
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11204 3896 11529 3924
rect 11204 3884 11210 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 11977 3927 12035 3933
rect 11977 3893 11989 3927
rect 12023 3924 12035 3927
rect 12526 3924 12532 3936
rect 12023 3896 12532 3924
rect 12023 3893 12035 3896
rect 11977 3887 12035 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 14182 3924 14188 3936
rect 14143 3896 14188 3924
rect 14182 3884 14188 3896
rect 14240 3884 14246 3936
rect 1104 3834 16468 3856
rect 1104 3782 3542 3834
rect 3594 3782 3606 3834
rect 3658 3782 3670 3834
rect 3722 3782 3734 3834
rect 3786 3782 8664 3834
rect 8716 3782 8728 3834
rect 8780 3782 8792 3834
rect 8844 3782 8856 3834
rect 8908 3782 13785 3834
rect 13837 3782 13849 3834
rect 13901 3782 13913 3834
rect 13965 3782 13977 3834
rect 14029 3782 16468 3834
rect 1104 3760 16468 3782
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 5215 3692 7052 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 3789 3655 3847 3661
rect 3789 3652 3801 3655
rect 2884 3624 3801 3652
rect 1946 3544 1952 3596
rect 2004 3584 2010 3596
rect 2041 3587 2099 3593
rect 2041 3584 2053 3587
rect 2004 3556 2053 3584
rect 2004 3544 2010 3556
rect 2041 3553 2053 3556
rect 2087 3553 2099 3587
rect 2041 3547 2099 3553
rect 2314 3544 2320 3596
rect 2372 3584 2378 3596
rect 2884 3593 2912 3624
rect 3789 3621 3801 3624
rect 3835 3621 3847 3655
rect 3789 3615 3847 3621
rect 4338 3612 4344 3664
rect 4396 3612 4402 3664
rect 4522 3612 4528 3664
rect 4580 3652 4586 3664
rect 5718 3652 5724 3664
rect 4580 3624 5724 3652
rect 4580 3612 4586 3624
rect 5718 3612 5724 3624
rect 5776 3652 5782 3664
rect 5902 3652 5908 3664
rect 5776 3624 5908 3652
rect 5776 3612 5782 3624
rect 5902 3612 5908 3624
rect 5960 3612 5966 3664
rect 7024 3652 7052 3692
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7653 3723 7711 3729
rect 7653 3720 7665 3723
rect 7156 3692 7665 3720
rect 7156 3680 7162 3692
rect 7653 3689 7665 3692
rect 7699 3689 7711 3723
rect 7653 3683 7711 3689
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 9122 3720 9128 3732
rect 8352 3692 9128 3720
rect 8352 3680 8358 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9490 3720 9496 3732
rect 9451 3692 9496 3720
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 10597 3723 10655 3729
rect 10597 3689 10609 3723
rect 10643 3720 10655 3723
rect 11149 3723 11207 3729
rect 11149 3720 11161 3723
rect 10643 3692 11161 3720
rect 10643 3689 10655 3692
rect 10597 3683 10655 3689
rect 11149 3689 11161 3692
rect 11195 3689 11207 3723
rect 11149 3683 11207 3689
rect 12802 3680 12808 3732
rect 12860 3720 12866 3732
rect 13538 3720 13544 3732
rect 12860 3692 13544 3720
rect 12860 3680 12866 3692
rect 13538 3680 13544 3692
rect 13596 3720 13602 3732
rect 14274 3720 14280 3732
rect 13596 3692 14280 3720
rect 13596 3680 13602 3692
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 15289 3723 15347 3729
rect 15289 3689 15301 3723
rect 15335 3720 15347 3723
rect 15378 3720 15384 3732
rect 15335 3692 15384 3720
rect 15335 3689 15347 3692
rect 15289 3683 15347 3689
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 8018 3652 8024 3664
rect 7024 3624 8024 3652
rect 8018 3612 8024 3624
rect 8076 3652 8082 3664
rect 8478 3652 8484 3664
rect 8076 3624 8156 3652
rect 8076 3612 8082 3624
rect 2409 3587 2467 3593
rect 2409 3584 2421 3587
rect 2372 3556 2421 3584
rect 2372 3544 2378 3556
rect 2409 3553 2421 3556
rect 2455 3553 2467 3587
rect 2409 3547 2467 3553
rect 2869 3587 2927 3593
rect 2869 3553 2881 3587
rect 2915 3553 2927 3587
rect 2869 3547 2927 3553
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 4356 3584 4384 3612
rect 8128 3593 8156 3624
rect 8312 3624 8484 3652
rect 8312 3593 8340 3624
rect 8478 3612 8484 3624
rect 8536 3652 8542 3664
rect 8536 3624 9674 3652
rect 8536 3612 8542 3624
rect 4433 3587 4491 3593
rect 4433 3584 4445 3587
rect 3200 3556 4108 3584
rect 4356 3556 4445 3584
rect 3200 3544 3206 3556
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 1854 3476 1860 3528
rect 1912 3516 1918 3528
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 1912 3488 2237 3516
rect 1912 3476 1918 3488
rect 2225 3485 2237 3488
rect 2271 3485 2283 3519
rect 2225 3479 2283 3485
rect 3878 3476 3884 3528
rect 3936 3525 3942 3528
rect 3936 3519 3972 3525
rect 3960 3485 3972 3519
rect 4080 3516 4108 3556
rect 4433 3553 4445 3556
rect 4479 3553 4491 3587
rect 8113 3587 8171 3593
rect 4433 3547 4491 3553
rect 5000 3556 7696 3584
rect 5000 3525 5028 3556
rect 4341 3519 4399 3525
rect 4341 3516 4353 3519
rect 4080 3488 4353 3516
rect 3936 3479 3972 3485
rect 4341 3485 4353 3488
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3485 5043 3519
rect 5166 3516 5172 3528
rect 5127 3488 5172 3516
rect 4985 3479 5043 3485
rect 3936 3476 3942 3479
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 5626 3476 5632 3528
rect 5684 3516 5690 3528
rect 5902 3516 5908 3528
rect 5684 3488 5729 3516
rect 5863 3488 5908 3516
rect 5684 3476 5690 3488
rect 5902 3476 5908 3488
rect 5960 3476 5966 3528
rect 5997 3519 6055 3525
rect 5997 3485 6009 3519
rect 6043 3516 6055 3519
rect 6086 3516 6092 3528
rect 6043 3488 6092 3516
rect 6043 3485 6055 3488
rect 5997 3479 6055 3485
rect 6086 3476 6092 3488
rect 6144 3476 6150 3528
rect 6730 3476 6736 3528
rect 6788 3516 6794 3528
rect 7009 3519 7067 3525
rect 7009 3516 7021 3519
rect 6788 3488 7021 3516
rect 6788 3476 6794 3488
rect 7009 3485 7021 3488
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 1489 3451 1547 3457
rect 1489 3417 1501 3451
rect 1535 3448 1547 3451
rect 5258 3448 5264 3460
rect 1535 3420 5264 3448
rect 1535 3417 1547 3420
rect 1489 3411 1547 3417
rect 5258 3408 5264 3420
rect 5316 3408 5322 3460
rect 5813 3451 5871 3457
rect 5813 3417 5825 3451
rect 5859 3417 5871 3451
rect 6822 3448 6828 3460
rect 6735 3420 6828 3448
rect 5813 3411 5871 3417
rect 2869 3383 2927 3389
rect 2869 3349 2881 3383
rect 2915 3380 2927 3383
rect 3510 3380 3516 3392
rect 2915 3352 3516 3380
rect 2915 3349 2927 3352
rect 2869 3343 2927 3349
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 3973 3383 4031 3389
rect 3973 3349 3985 3383
rect 4019 3380 4031 3383
rect 4062 3380 4068 3392
rect 4019 3352 4068 3380
rect 4019 3349 4031 3352
rect 3973 3343 4031 3349
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 5442 3340 5448 3392
rect 5500 3380 5506 3392
rect 5828 3380 5856 3411
rect 6822 3408 6828 3420
rect 6880 3448 6886 3460
rect 7190 3448 7196 3460
rect 6880 3420 7196 3448
rect 6880 3408 6886 3420
rect 7190 3408 7196 3420
rect 7248 3408 7254 3460
rect 7668 3448 7696 3556
rect 8113 3553 8125 3587
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 8297 3587 8355 3593
rect 8297 3553 8309 3587
rect 8343 3553 8355 3587
rect 8297 3547 8355 3553
rect 9033 3587 9091 3593
rect 9033 3553 9045 3587
rect 9079 3584 9091 3587
rect 9398 3584 9404 3596
rect 9079 3556 9404 3584
rect 9079 3553 9091 3556
rect 9033 3547 9091 3553
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 9646 3584 9674 3624
rect 10318 3612 10324 3664
rect 10376 3652 10382 3664
rect 11609 3655 11667 3661
rect 11609 3652 11621 3655
rect 10376 3624 11621 3652
rect 10376 3612 10382 3624
rect 11609 3621 11621 3624
rect 11655 3652 11667 3655
rect 11790 3652 11796 3664
rect 11655 3624 11796 3652
rect 11655 3621 11667 3624
rect 11609 3615 11667 3621
rect 11790 3612 11796 3624
rect 11848 3612 11854 3664
rect 12618 3612 12624 3664
rect 12676 3652 12682 3664
rect 12897 3655 12955 3661
rect 12897 3652 12909 3655
rect 12676 3624 12909 3652
rect 12676 3612 12682 3624
rect 12897 3621 12909 3624
rect 12943 3621 12955 3655
rect 12897 3615 12955 3621
rect 13357 3655 13415 3661
rect 13357 3621 13369 3655
rect 13403 3652 13415 3655
rect 13403 3624 14780 3652
rect 13403 3621 13415 3624
rect 13357 3615 13415 3621
rect 11514 3584 11520 3596
rect 9646 3556 10732 3584
rect 11427 3556 11520 3584
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8662 3516 8668 3528
rect 8260 3488 8668 3516
rect 8260 3476 8266 3488
rect 8662 3476 8668 3488
rect 8720 3516 8726 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8720 3488 8953 3516
rect 8720 3476 8726 3488
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 9214 3516 9220 3528
rect 9175 3488 9220 3516
rect 8941 3479 8999 3485
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 10704 3525 10732 3556
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 10689 3519 10747 3525
rect 10689 3485 10701 3519
rect 10735 3516 10747 3519
rect 11146 3516 11152 3528
rect 10735 3488 11152 3516
rect 10735 3485 10747 3488
rect 10689 3479 10747 3485
rect 9324 3448 9352 3479
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 11440 3525 11468 3556
rect 11514 3544 11520 3556
rect 11572 3584 11578 3596
rect 12158 3584 12164 3596
rect 11572 3556 12164 3584
rect 11572 3544 11578 3556
rect 12158 3544 12164 3556
rect 12216 3544 12222 3596
rect 14182 3584 14188 3596
rect 12452 3556 14188 3584
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3485 11391 3519
rect 11333 3479 11391 3485
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3485 11483 3519
rect 11425 3479 11483 3485
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3516 11759 3519
rect 12342 3516 12348 3528
rect 11747 3488 12348 3516
rect 11747 3485 11759 3488
rect 11701 3479 11759 3485
rect 11348 3448 11376 3479
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 12452 3525 12480 3556
rect 13464 3525 13492 3556
rect 14182 3544 14188 3556
rect 14240 3584 14246 3596
rect 14752 3593 14780 3624
rect 14737 3587 14795 3593
rect 14240 3556 14504 3584
rect 14240 3544 14246 3556
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3485 12495 3519
rect 12437 3479 12495 3485
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3485 13231 3519
rect 13173 3479 13231 3485
rect 13449 3519 13507 3525
rect 13449 3485 13461 3519
rect 13495 3485 13507 3519
rect 13449 3479 13507 3485
rect 12710 3448 12716 3460
rect 7668 3420 12716 3448
rect 12710 3408 12716 3420
rect 12768 3408 12774 3460
rect 5500 3352 5856 3380
rect 5500 3340 5506 3352
rect 5994 3340 6000 3392
rect 6052 3380 6058 3392
rect 6181 3383 6239 3389
rect 6181 3380 6193 3383
rect 6052 3352 6193 3380
rect 6052 3340 6058 3352
rect 6181 3349 6193 3352
rect 6227 3349 6239 3383
rect 6181 3343 6239 3349
rect 6546 3340 6552 3392
rect 6604 3380 6610 3392
rect 6641 3383 6699 3389
rect 6641 3380 6653 3383
rect 6604 3352 6653 3380
rect 6604 3340 6610 3352
rect 6641 3349 6653 3352
rect 6687 3349 6699 3383
rect 6641 3343 6699 3349
rect 8021 3383 8079 3389
rect 8021 3349 8033 3383
rect 8067 3380 8079 3383
rect 8386 3380 8392 3392
rect 8067 3352 8392 3380
rect 8067 3349 8079 3352
rect 8021 3343 8079 3349
rect 8386 3340 8392 3352
rect 8444 3340 8450 3392
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 10229 3383 10287 3389
rect 10229 3380 10241 3383
rect 9364 3352 10241 3380
rect 9364 3340 9370 3352
rect 10229 3349 10241 3352
rect 10275 3349 10287 3383
rect 10229 3343 10287 3349
rect 12345 3383 12403 3389
rect 12345 3349 12357 3383
rect 12391 3380 12403 3383
rect 12802 3380 12808 3392
rect 12391 3352 12808 3380
rect 12391 3349 12403 3352
rect 12345 3343 12403 3349
rect 12802 3340 12808 3352
rect 12860 3340 12866 3392
rect 13096 3380 13124 3479
rect 13188 3448 13216 3479
rect 14274 3476 14280 3528
rect 14332 3516 14338 3528
rect 14476 3516 14504 3556
rect 14737 3553 14749 3587
rect 14783 3584 14795 3587
rect 14826 3584 14832 3596
rect 14783 3556 14832 3584
rect 14783 3553 14795 3556
rect 14737 3547 14795 3553
rect 14826 3544 14832 3556
rect 14884 3544 14890 3596
rect 14579 3519 14637 3525
rect 14579 3516 14591 3519
rect 14332 3488 14377 3516
rect 14476 3488 14591 3516
rect 14332 3476 14338 3488
rect 14579 3485 14591 3488
rect 14625 3485 14637 3519
rect 14579 3479 14637 3485
rect 15102 3476 15108 3528
rect 15160 3516 15166 3528
rect 15197 3519 15255 3525
rect 15197 3516 15209 3519
rect 15160 3488 15209 3516
rect 15160 3476 15166 3488
rect 15197 3485 15209 3488
rect 15243 3485 15255 3519
rect 15197 3479 15255 3485
rect 14369 3451 14427 3457
rect 13188 3420 13952 3448
rect 13924 3392 13952 3420
rect 14369 3417 14381 3451
rect 14415 3417 14427 3451
rect 14369 3411 14427 3417
rect 13814 3380 13820 3392
rect 13096 3352 13820 3380
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 13906 3340 13912 3392
rect 13964 3380 13970 3392
rect 14093 3383 14151 3389
rect 14093 3380 14105 3383
rect 13964 3352 14105 3380
rect 13964 3340 13970 3352
rect 14093 3349 14105 3352
rect 14139 3349 14151 3383
rect 14384 3380 14412 3411
rect 14458 3408 14464 3460
rect 14516 3448 14522 3460
rect 14516 3420 14561 3448
rect 14516 3408 14522 3420
rect 14918 3380 14924 3392
rect 14384 3352 14924 3380
rect 14093 3343 14151 3349
rect 14918 3340 14924 3352
rect 14976 3340 14982 3392
rect 1104 3290 16468 3312
rect 1104 3238 6103 3290
rect 6155 3238 6167 3290
rect 6219 3238 6231 3290
rect 6283 3238 6295 3290
rect 6347 3238 11224 3290
rect 11276 3238 11288 3290
rect 11340 3238 11352 3290
rect 11404 3238 11416 3290
rect 11468 3238 16468 3290
rect 1104 3216 16468 3238
rect 2590 3176 2596 3188
rect 2551 3148 2596 3176
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 4062 3136 4068 3188
rect 4120 3136 4126 3188
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 5316 3148 8432 3176
rect 5316 3136 5322 3148
rect 1394 3108 1400 3120
rect 1355 3080 1400 3108
rect 1394 3068 1400 3080
rect 1452 3108 1458 3120
rect 3326 3108 3332 3120
rect 1452 3080 1900 3108
rect 3287 3080 3332 3108
rect 1452 3068 1458 3080
rect 1489 3043 1547 3049
rect 1489 3009 1501 3043
rect 1535 3040 1547 3043
rect 1762 3040 1768 3052
rect 1535 3012 1768 3040
rect 1535 3009 1547 3012
rect 1489 3003 1547 3009
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 1872 3049 1900 3080
rect 3326 3068 3332 3080
rect 3384 3068 3390 3120
rect 4080 3108 4108 3136
rect 3436 3080 4108 3108
rect 4341 3111 4399 3117
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2682 3000 2688 3052
rect 2740 3038 2746 3052
rect 3142 3040 3148 3052
rect 2740 3010 2783 3038
rect 3055 3012 3148 3040
rect 2740 3000 2746 3010
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 3436 3049 3464 3080
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 7282 3108 7288 3120
rect 4387 3080 7288 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 3510 3000 3516 3052
rect 3568 3040 3574 3052
rect 4065 3043 4123 3049
rect 4065 3040 4077 3043
rect 3568 3012 4077 3040
rect 3568 3000 3574 3012
rect 4065 3009 4077 3012
rect 4111 3040 4123 3043
rect 4356 3040 4384 3071
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 4111 3012 4384 3040
rect 5445 3043 5503 3049
rect 4111 3009 4123 3012
rect 4065 3003 4123 3009
rect 5445 3009 5457 3043
rect 5491 3040 5503 3043
rect 5721 3043 5779 3049
rect 5721 3040 5733 3043
rect 5491 3012 5733 3040
rect 5491 3009 5503 3012
rect 5445 3003 5503 3009
rect 2130 2932 2136 2984
rect 2188 2972 2194 2984
rect 3160 2972 3188 3000
rect 5552 2984 5580 3012
rect 5721 3009 5733 3012
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 7193 3043 7251 3049
rect 7193 3040 7205 3043
rect 5960 3012 7205 3040
rect 5960 3000 5966 3012
rect 7193 3009 7205 3012
rect 7239 3040 7251 3043
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 7239 3012 7481 3040
rect 7239 3009 7251 3012
rect 7193 3003 7251 3009
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 8404 3049 8432 3148
rect 9122 3136 9128 3188
rect 9180 3176 9186 3188
rect 11514 3176 11520 3188
rect 9180 3148 11520 3176
rect 9180 3136 9186 3148
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 11701 3179 11759 3185
rect 11701 3145 11713 3179
rect 11747 3176 11759 3179
rect 11747 3148 12434 3176
rect 11747 3145 11759 3148
rect 11701 3139 11759 3145
rect 8754 3068 8760 3120
rect 8812 3108 8818 3120
rect 12406 3108 12434 3148
rect 13170 3136 13176 3188
rect 13228 3176 13234 3188
rect 17494 3176 17500 3188
rect 13228 3148 17500 3176
rect 13228 3136 13234 3148
rect 17494 3136 17500 3148
rect 17552 3136 17558 3188
rect 12526 3108 12532 3120
rect 8812 3080 10180 3108
rect 12406 3080 12532 3108
rect 8812 3068 8818 3080
rect 8205 3043 8263 3049
rect 8205 3040 8217 3043
rect 7892 3012 8217 3040
rect 7892 3000 7898 3012
rect 8205 3009 8217 3012
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 8536 3012 8581 3040
rect 8536 3000 8542 3012
rect 8662 3000 8668 3052
rect 8720 3040 8726 3052
rect 9674 3040 9680 3052
rect 8720 3012 8765 3040
rect 9635 3012 9680 3040
rect 8720 3000 8726 3012
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 10152 3049 10180 3080
rect 12526 3068 12532 3080
rect 12584 3108 12590 3120
rect 12802 3108 12808 3120
rect 12584 3080 12808 3108
rect 12584 3068 12590 3080
rect 12802 3068 12808 3080
rect 12860 3108 12866 3120
rect 13446 3108 13452 3120
rect 12860 3080 13452 3108
rect 12860 3068 12866 3080
rect 13446 3068 13452 3080
rect 13504 3068 13510 3120
rect 13538 3068 13544 3120
rect 13596 3068 13602 3120
rect 13906 3108 13912 3120
rect 13648 3080 13912 3108
rect 10137 3043 10195 3049
rect 10137 3009 10149 3043
rect 10183 3009 10195 3043
rect 10502 3040 10508 3052
rect 10463 3012 10508 3040
rect 10137 3003 10195 3009
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11112 3012 11529 3040
rect 11112 3000 11118 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 12250 3040 12256 3052
rect 12211 3012 12256 3040
rect 11517 3003 11575 3009
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 13262 3000 13268 3052
rect 13320 3040 13326 3052
rect 13556 3040 13584 3068
rect 13648 3049 13676 3080
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 14001 3111 14059 3117
rect 14001 3077 14013 3111
rect 14047 3108 14059 3111
rect 14090 3108 14096 3120
rect 14047 3080 14096 3108
rect 14047 3077 14059 3080
rect 14001 3071 14059 3077
rect 13320 3012 13584 3040
rect 13633 3043 13691 3049
rect 13320 3000 13326 3012
rect 13633 3009 13645 3043
rect 13679 3009 13691 3043
rect 13633 3003 13691 3009
rect 2188 2944 3188 2972
rect 3881 2975 3939 2981
rect 2188 2932 2194 2944
rect 3881 2941 3893 2975
rect 3927 2972 3939 2975
rect 4430 2972 4436 2984
rect 3927 2944 4436 2972
rect 3927 2941 3939 2944
rect 3881 2935 3939 2941
rect 4430 2932 4436 2944
rect 4488 2932 4494 2984
rect 5353 2975 5411 2981
rect 5353 2941 5365 2975
rect 5399 2941 5411 2975
rect 5353 2935 5411 2941
rect 2041 2907 2099 2913
rect 2041 2873 2053 2907
rect 2087 2904 2099 2907
rect 4062 2904 4068 2916
rect 2087 2876 4068 2904
rect 2087 2873 2099 2876
rect 2041 2867 2099 2873
rect 4062 2864 4068 2876
rect 4120 2864 4126 2916
rect 4157 2907 4215 2913
rect 4157 2873 4169 2907
rect 4203 2904 4215 2907
rect 4246 2904 4252 2916
rect 4203 2876 4252 2904
rect 4203 2873 4215 2876
rect 4157 2867 4215 2873
rect 4246 2864 4252 2876
rect 4304 2864 4310 2916
rect 5368 2904 5396 2935
rect 5534 2932 5540 2984
rect 5592 2932 5598 2984
rect 5813 2975 5871 2981
rect 5813 2941 5825 2975
rect 5859 2972 5871 2975
rect 5994 2972 6000 2984
rect 5859 2944 6000 2972
rect 5859 2941 5871 2944
rect 5813 2935 5871 2941
rect 5828 2904 5856 2935
rect 5994 2932 6000 2944
rect 6052 2972 6058 2984
rect 6730 2972 6736 2984
rect 6052 2944 6736 2972
rect 6052 2932 6058 2944
rect 6730 2932 6736 2944
rect 6788 2932 6794 2984
rect 6822 2932 6828 2984
rect 6880 2932 6886 2984
rect 7098 2972 7104 2984
rect 7059 2944 7104 2972
rect 7098 2932 7104 2944
rect 7156 2972 7162 2984
rect 7561 2975 7619 2981
rect 7561 2972 7573 2975
rect 7156 2944 7573 2972
rect 7156 2932 7162 2944
rect 7561 2941 7573 2944
rect 7607 2941 7619 2975
rect 9858 2972 9864 2984
rect 7561 2935 7619 2941
rect 7668 2944 9864 2972
rect 5368 2876 5856 2904
rect 1854 2796 1860 2848
rect 1912 2836 1918 2848
rect 3145 2839 3203 2845
rect 3145 2836 3157 2839
rect 1912 2808 3157 2836
rect 1912 2796 1918 2808
rect 3145 2805 3157 2808
rect 3191 2805 3203 2839
rect 3145 2799 3203 2805
rect 3878 2796 3884 2848
rect 3936 2836 3942 2848
rect 5169 2839 5227 2845
rect 5169 2836 5181 2839
rect 3936 2808 5181 2836
rect 3936 2796 3942 2808
rect 5169 2805 5181 2808
rect 5215 2805 5227 2839
rect 6849 2836 6877 2932
rect 7006 2864 7012 2916
rect 7064 2904 7070 2916
rect 7668 2904 7696 2944
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 9950 2932 9956 2984
rect 10008 2972 10014 2984
rect 10413 2975 10471 2981
rect 10413 2972 10425 2975
rect 10008 2944 10425 2972
rect 10008 2932 10014 2944
rect 10413 2941 10425 2944
rect 10459 2941 10471 2975
rect 10413 2935 10471 2941
rect 12805 2975 12863 2981
rect 12805 2941 12817 2975
rect 12851 2972 12863 2975
rect 12894 2972 12900 2984
rect 12851 2944 12900 2972
rect 12851 2941 12863 2944
rect 12805 2935 12863 2941
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 13541 2975 13599 2981
rect 13541 2941 13553 2975
rect 13587 2972 13599 2975
rect 13814 2972 13820 2984
rect 13587 2944 13820 2972
rect 13587 2941 13599 2944
rect 13541 2935 13599 2941
rect 13814 2932 13820 2944
rect 13872 2972 13878 2984
rect 14016 2972 14044 3071
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 14826 3108 14832 3120
rect 14200 3080 14596 3108
rect 14787 3080 14832 3108
rect 13872 2944 14044 2972
rect 13872 2932 13878 2944
rect 7064 2876 7696 2904
rect 7064 2864 7070 2876
rect 7742 2864 7748 2916
rect 7800 2904 7806 2916
rect 8297 2907 8355 2913
rect 7800 2876 8248 2904
rect 7800 2864 7806 2876
rect 6917 2839 6975 2845
rect 6917 2836 6929 2839
rect 6849 2808 6929 2836
rect 5169 2799 5227 2805
rect 6917 2805 6929 2808
rect 6963 2805 6975 2839
rect 6917 2799 6975 2805
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 8021 2839 8079 2845
rect 8021 2836 8033 2839
rect 7156 2808 8033 2836
rect 7156 2796 7162 2808
rect 8021 2805 8033 2808
rect 8067 2805 8079 2839
rect 8220 2836 8248 2876
rect 8297 2873 8309 2907
rect 8343 2904 8355 2907
rect 8386 2904 8392 2916
rect 8343 2876 8392 2904
rect 8343 2873 8355 2876
rect 8297 2867 8355 2873
rect 8386 2864 8392 2876
rect 8444 2904 8450 2916
rect 9214 2904 9220 2916
rect 8444 2876 9220 2904
rect 8444 2864 8450 2876
rect 9214 2864 9220 2876
rect 9272 2864 9278 2916
rect 10321 2907 10379 2913
rect 10321 2873 10333 2907
rect 10367 2904 10379 2907
rect 14200 2904 14228 3080
rect 14461 3043 14519 3049
rect 14461 3009 14473 3043
rect 14507 3009 14519 3043
rect 14461 3003 14519 3009
rect 10367 2876 14228 2904
rect 10367 2873 10379 2876
rect 10321 2867 10379 2873
rect 13170 2836 13176 2848
rect 8220 2808 13176 2836
rect 8021 2799 8079 2805
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 13262 2796 13268 2848
rect 13320 2836 13326 2848
rect 13357 2839 13415 2845
rect 13357 2836 13369 2839
rect 13320 2808 13369 2836
rect 13320 2796 13326 2808
rect 13357 2805 13369 2808
rect 13403 2805 13415 2839
rect 13357 2799 13415 2805
rect 13446 2796 13452 2848
rect 13504 2836 13510 2848
rect 14476 2836 14504 3003
rect 14568 2972 14596 3080
rect 14826 3068 14832 3080
rect 14884 3068 14890 3120
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3040 14703 3043
rect 15378 3040 15384 3052
rect 14691 3012 15384 3040
rect 14691 3009 14703 3012
rect 14645 3003 14703 3009
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 15565 3043 15623 3049
rect 15565 3009 15577 3043
rect 15611 3009 15623 3043
rect 15565 3003 15623 3009
rect 15580 2972 15608 3003
rect 14568 2944 15608 2972
rect 15746 2904 15752 2916
rect 15707 2876 15752 2904
rect 15746 2864 15752 2876
rect 15804 2864 15810 2916
rect 13504 2808 14504 2836
rect 13504 2796 13510 2808
rect 1104 2746 16468 2768
rect 1104 2694 3542 2746
rect 3594 2694 3606 2746
rect 3658 2694 3670 2746
rect 3722 2694 3734 2746
rect 3786 2694 8664 2746
rect 8716 2694 8728 2746
rect 8780 2694 8792 2746
rect 8844 2694 8856 2746
rect 8908 2694 13785 2746
rect 13837 2694 13849 2746
rect 13901 2694 13913 2746
rect 13965 2694 13977 2746
rect 14029 2694 16468 2746
rect 1104 2672 16468 2694
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5902 2632 5908 2644
rect 4939 2604 5908 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 5902 2592 5908 2604
rect 5960 2592 5966 2644
rect 6457 2635 6515 2641
rect 6457 2601 6469 2635
rect 6503 2632 6515 2635
rect 6914 2632 6920 2644
rect 6503 2604 6920 2632
rect 6503 2601 6515 2604
rect 6457 2595 6515 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7466 2632 7472 2644
rect 7427 2604 7472 2632
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 8205 2635 8263 2641
rect 8205 2601 8217 2635
rect 8251 2601 8263 2635
rect 8205 2595 8263 2601
rect 4706 2524 4712 2576
rect 4764 2564 4770 2576
rect 8220 2564 8248 2595
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8352 2604 8953 2632
rect 8352 2592 8358 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 9858 2632 9864 2644
rect 9815 2604 9864 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 11790 2632 11796 2644
rect 9968 2604 11796 2632
rect 8389 2567 8447 2573
rect 4764 2536 8340 2564
rect 4764 2524 4770 2536
rect 2038 2456 2044 2508
rect 2096 2496 2102 2508
rect 4798 2496 4804 2508
rect 2096 2468 4804 2496
rect 2096 2456 2102 2468
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1397 2391 1455 2397
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 2958 2428 2964 2440
rect 2915 2400 2964 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 4908 2437 4936 2536
rect 8312 2508 8340 2536
rect 8389 2533 8401 2567
rect 8435 2533 8447 2567
rect 8389 2527 8447 2533
rect 5626 2456 5632 2508
rect 5684 2496 5690 2508
rect 6546 2496 6552 2508
rect 5684 2468 6552 2496
rect 5684 2456 5690 2468
rect 4341 2431 4399 2437
rect 4341 2428 4353 2431
rect 4120 2400 4353 2428
rect 4120 2388 4126 2400
rect 4341 2397 4353 2400
rect 4387 2397 4399 2431
rect 4341 2391 4399 2397
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 5442 2428 5448 2440
rect 5123 2400 5448 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2428 5779 2431
rect 5810 2428 5816 2440
rect 5767 2400 5816 2428
rect 5767 2397 5779 2400
rect 5721 2391 5779 2397
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6380 2437 6408 2468
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 8294 2456 8300 2508
rect 8352 2456 8358 2508
rect 8404 2496 8432 2527
rect 9398 2524 9404 2576
rect 9456 2564 9462 2576
rect 9968 2564 9996 2604
rect 11790 2592 11796 2604
rect 11848 2632 11854 2644
rect 12621 2635 12679 2641
rect 12621 2632 12633 2635
rect 11848 2604 12633 2632
rect 11848 2592 11854 2604
rect 12621 2601 12633 2604
rect 12667 2601 12679 2635
rect 12621 2595 12679 2601
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 13265 2635 13323 2641
rect 13265 2632 13277 2635
rect 12768 2604 13277 2632
rect 12768 2592 12774 2604
rect 13265 2601 13277 2604
rect 13311 2601 13323 2635
rect 13265 2595 13323 2601
rect 13909 2635 13967 2641
rect 13909 2601 13921 2635
rect 13955 2632 13967 2635
rect 14185 2635 14243 2641
rect 14185 2632 14197 2635
rect 13955 2604 14197 2632
rect 13955 2601 13967 2604
rect 13909 2595 13967 2601
rect 14185 2601 14197 2604
rect 14231 2632 14243 2635
rect 14642 2632 14648 2644
rect 14231 2604 14648 2632
rect 14231 2601 14243 2604
rect 14185 2595 14243 2601
rect 14642 2592 14648 2604
rect 14700 2592 14706 2644
rect 9456 2536 9996 2564
rect 9456 2524 9462 2536
rect 10042 2524 10048 2576
rect 10100 2564 10106 2576
rect 10100 2536 12112 2564
rect 10100 2524 10106 2536
rect 10321 2499 10379 2505
rect 10321 2496 10333 2499
rect 8404 2468 10333 2496
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 6641 2431 6699 2437
rect 6641 2422 6653 2431
rect 6365 2391 6423 2397
rect 6564 2397 6653 2422
rect 6687 2397 6699 2431
rect 6564 2394 6699 2397
rect 1854 2320 1860 2372
rect 1912 2360 1918 2372
rect 2685 2363 2743 2369
rect 2685 2360 2697 2363
rect 1912 2332 2697 2360
rect 1912 2320 1918 2332
rect 2685 2329 2697 2332
rect 2731 2329 2743 2363
rect 2685 2323 2743 2329
rect 3878 2320 3884 2372
rect 3936 2360 3942 2372
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 3936 2332 4169 2360
rect 3936 2320 3942 2332
rect 4157 2329 4169 2332
rect 4203 2329 4215 2363
rect 4157 2323 4215 2329
rect 5534 2320 5540 2372
rect 5592 2360 5598 2372
rect 6564 2360 6592 2394
rect 6641 2391 6699 2394
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 7558 2428 7564 2440
rect 6788 2400 6833 2428
rect 7519 2400 7564 2428
rect 6788 2388 6794 2400
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 8018 2428 8024 2440
rect 7979 2400 8024 2428
rect 8018 2388 8024 2400
rect 8076 2388 8082 2440
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 9122 2428 9128 2440
rect 9083 2400 9128 2428
rect 8205 2391 8263 2397
rect 7098 2360 7104 2372
rect 5592 2332 7104 2360
rect 5592 2320 5598 2332
rect 7098 2320 7104 2332
rect 7156 2320 7162 2372
rect 8220 2360 8248 2391
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 9950 2428 9956 2440
rect 9508 2400 9956 2428
rect 9309 2363 9367 2369
rect 9309 2360 9321 2363
rect 8220 2332 9321 2360
rect 9309 2329 9321 2332
rect 9355 2360 9367 2363
rect 9398 2360 9404 2372
rect 9355 2332 9404 2360
rect 9355 2329 9367 2332
rect 9309 2323 9367 2329
rect 9398 2320 9404 2332
rect 9456 2320 9462 2372
rect 5626 2292 5632 2304
rect 5587 2264 5632 2292
rect 5626 2252 5632 2264
rect 5684 2252 5690 2304
rect 6917 2295 6975 2301
rect 6917 2261 6929 2295
rect 6963 2292 6975 2295
rect 9508 2292 9536 2400
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 10060 2437 10088 2468
rect 10321 2465 10333 2468
rect 10367 2496 10379 2499
rect 10502 2496 10508 2508
rect 10367 2468 10508 2496
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 10502 2456 10508 2468
rect 10560 2456 10566 2508
rect 12084 2437 12112 2536
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14384 2468 14933 2496
rect 14384 2440 14412 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2397 10103 2431
rect 10045 2391 10103 2397
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2397 12127 2431
rect 12802 2428 12808 2440
rect 12763 2400 12808 2428
rect 12069 2391 12127 2397
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2428 13507 2431
rect 13909 2431 13967 2437
rect 13909 2428 13921 2431
rect 13495 2400 13921 2428
rect 13495 2397 13507 2400
rect 13449 2391 13507 2397
rect 13909 2397 13921 2400
rect 13955 2397 13967 2431
rect 14366 2428 14372 2440
rect 14327 2400 14372 2428
rect 13909 2391 13967 2397
rect 14366 2388 14372 2400
rect 14424 2388 14430 2440
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 9968 2360 9996 2388
rect 10413 2363 10471 2369
rect 10413 2360 10425 2363
rect 9968 2332 10425 2360
rect 10413 2329 10425 2332
rect 10459 2329 10471 2363
rect 10413 2323 10471 2329
rect 13354 2320 13360 2372
rect 13412 2360 13418 2372
rect 14844 2360 14872 2391
rect 15470 2360 15476 2372
rect 13412 2332 14872 2360
rect 15431 2332 15476 2360
rect 13412 2320 13418 2332
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 15654 2360 15660 2372
rect 15615 2332 15660 2360
rect 15654 2320 15660 2332
rect 15712 2320 15718 2372
rect 6963 2264 9536 2292
rect 6963 2261 6975 2264
rect 6917 2255 6975 2261
rect 9582 2252 9588 2304
rect 9640 2292 9646 2304
rect 11977 2295 12035 2301
rect 11977 2292 11989 2295
rect 9640 2264 11989 2292
rect 9640 2252 9646 2264
rect 11977 2261 11989 2264
rect 12023 2261 12035 2295
rect 11977 2255 12035 2261
rect 1104 2202 16468 2224
rect 1104 2150 6103 2202
rect 6155 2150 6167 2202
rect 6219 2150 6231 2202
rect 6283 2150 6295 2202
rect 6347 2150 11224 2202
rect 11276 2150 11288 2202
rect 11340 2150 11352 2202
rect 11404 2150 11416 2202
rect 11468 2150 16468 2202
rect 1104 2128 16468 2150
rect 1670 2048 1676 2100
rect 1728 2088 1734 2100
rect 9490 2088 9496 2100
rect 1728 2060 9496 2088
rect 1728 2048 1734 2060
rect 9490 2048 9496 2060
rect 9548 2048 9554 2100
rect 4798 1980 4804 2032
rect 4856 2020 4862 2032
rect 15654 2020 15660 2032
rect 4856 1992 15660 2020
rect 4856 1980 4862 1992
rect 15654 1980 15660 1992
rect 15712 1980 15718 2032
<< via1 >>
rect 6103 17382 6155 17434
rect 6167 17382 6219 17434
rect 6231 17382 6283 17434
rect 6295 17382 6347 17434
rect 11224 17382 11276 17434
rect 11288 17382 11340 17434
rect 11352 17382 11404 17434
rect 11416 17382 11468 17434
rect 20 17280 72 17332
rect 9772 17280 9824 17332
rect 1860 17255 1912 17264
rect 1860 17221 1869 17255
rect 1869 17221 1903 17255
rect 1903 17221 1912 17255
rect 1860 17212 1912 17221
rect 4160 17255 4212 17264
rect 4160 17221 4169 17255
rect 4169 17221 4203 17255
rect 4203 17221 4212 17255
rect 4160 17212 4212 17221
rect 7932 17212 7984 17264
rect 8300 17212 8352 17264
rect 11888 17212 11940 17264
rect 1676 17144 1728 17196
rect 4252 17144 4304 17196
rect 5080 17187 5132 17196
rect 5080 17153 5089 17187
rect 5089 17153 5123 17187
rect 5123 17153 5132 17187
rect 5080 17144 5132 17153
rect 5448 17144 5500 17196
rect 5908 17144 5960 17196
rect 8208 17187 8260 17196
rect 8208 17153 8217 17187
rect 8217 17153 8251 17187
rect 8251 17153 8260 17187
rect 8208 17144 8260 17153
rect 9404 17187 9456 17196
rect 4896 17051 4948 17060
rect 4896 17017 4905 17051
rect 4905 17017 4939 17051
rect 4939 17017 4948 17051
rect 4896 17008 4948 17017
rect 6920 17076 6972 17128
rect 9404 17153 9413 17187
rect 9413 17153 9447 17187
rect 9447 17153 9456 17187
rect 9404 17144 9456 17153
rect 10324 17144 10376 17196
rect 11704 17187 11756 17196
rect 9312 17076 9364 17128
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 11796 17187 11848 17196
rect 11796 17153 11805 17187
rect 11805 17153 11839 17187
rect 11839 17153 11848 17187
rect 12072 17187 12124 17196
rect 11796 17144 11848 17153
rect 12072 17153 12081 17187
rect 12081 17153 12115 17187
rect 12115 17153 12124 17187
rect 12072 17144 12124 17153
rect 12164 17144 12216 17196
rect 13820 17144 13872 17196
rect 17500 17212 17552 17264
rect 15384 17144 15436 17196
rect 7472 17008 7524 17060
rect 12900 17008 12952 17060
rect 15752 17051 15804 17060
rect 15752 17017 15761 17051
rect 15761 17017 15795 17051
rect 15795 17017 15804 17051
rect 15752 17008 15804 17017
rect 6092 16940 6144 16992
rect 8116 16940 8168 16992
rect 10232 16940 10284 16992
rect 11520 16983 11572 16992
rect 11520 16949 11529 16983
rect 11529 16949 11563 16983
rect 11563 16949 11572 16983
rect 11520 16940 11572 16949
rect 11888 16940 11940 16992
rect 12716 16940 12768 16992
rect 14556 16940 14608 16992
rect 3542 16838 3594 16890
rect 3606 16838 3658 16890
rect 3670 16838 3722 16890
rect 3734 16838 3786 16890
rect 8664 16838 8716 16890
rect 8728 16838 8780 16890
rect 8792 16838 8844 16890
rect 8856 16838 8908 16890
rect 13785 16838 13837 16890
rect 13849 16838 13901 16890
rect 13913 16838 13965 16890
rect 13977 16838 14029 16890
rect 5080 16736 5132 16788
rect 8208 16736 8260 16788
rect 11796 16736 11848 16788
rect 3056 16668 3108 16720
rect 2504 16532 2556 16584
rect 3700 16600 3752 16652
rect 7104 16600 7156 16652
rect 2780 16532 2832 16584
rect 4068 16532 4120 16584
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 4988 16532 5040 16541
rect 5356 16575 5408 16584
rect 5356 16541 5365 16575
rect 5365 16541 5399 16575
rect 5399 16541 5408 16575
rect 5356 16532 5408 16541
rect 5816 16575 5868 16584
rect 5816 16541 5825 16575
rect 5825 16541 5859 16575
rect 5859 16541 5868 16575
rect 5816 16532 5868 16541
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 7012 16575 7064 16584
rect 7012 16541 7021 16575
rect 7021 16541 7055 16575
rect 7055 16541 7064 16575
rect 7012 16532 7064 16541
rect 8300 16532 8352 16584
rect 8392 16575 8444 16584
rect 8392 16541 8401 16575
rect 8401 16541 8435 16575
rect 8435 16541 8444 16575
rect 9404 16575 9456 16584
rect 8392 16532 8444 16541
rect 9404 16541 9413 16575
rect 9413 16541 9447 16575
rect 9447 16541 9456 16575
rect 10416 16600 10468 16652
rect 12072 16600 12124 16652
rect 13452 16668 13504 16720
rect 13544 16643 13596 16652
rect 13544 16609 13553 16643
rect 13553 16609 13587 16643
rect 13587 16609 13596 16643
rect 13544 16600 13596 16609
rect 9404 16532 9456 16541
rect 10232 16575 10284 16584
rect 10232 16541 10241 16575
rect 10241 16541 10275 16575
rect 10275 16541 10284 16575
rect 10232 16532 10284 16541
rect 11888 16575 11940 16584
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 11888 16532 11940 16541
rect 14372 16575 14424 16584
rect 2044 16464 2096 16516
rect 4896 16464 4948 16516
rect 9220 16507 9272 16516
rect 2504 16439 2556 16448
rect 2504 16405 2513 16439
rect 2513 16405 2547 16439
rect 2547 16405 2556 16439
rect 2504 16396 2556 16405
rect 5448 16396 5500 16448
rect 5632 16396 5684 16448
rect 7564 16439 7616 16448
rect 7564 16405 7573 16439
rect 7573 16405 7607 16439
rect 7607 16405 7616 16439
rect 7564 16396 7616 16405
rect 8300 16439 8352 16448
rect 8300 16405 8309 16439
rect 8309 16405 8343 16439
rect 8343 16405 8352 16439
rect 8300 16396 8352 16405
rect 9220 16473 9229 16507
rect 9229 16473 9263 16507
rect 9263 16473 9272 16507
rect 9220 16464 9272 16473
rect 11520 16464 11572 16516
rect 14372 16541 14381 16575
rect 14381 16541 14415 16575
rect 14415 16541 14424 16575
rect 14372 16532 14424 16541
rect 14464 16575 14516 16584
rect 14464 16541 14473 16575
rect 14473 16541 14507 16575
rect 14507 16541 14516 16575
rect 14464 16532 14516 16541
rect 13452 16507 13504 16516
rect 13452 16473 13461 16507
rect 13461 16473 13495 16507
rect 13495 16473 13504 16507
rect 13452 16464 13504 16473
rect 15200 16507 15252 16516
rect 15200 16473 15209 16507
rect 15209 16473 15243 16507
rect 15243 16473 15252 16507
rect 15200 16464 15252 16473
rect 15292 16464 15344 16516
rect 12164 16396 12216 16448
rect 14372 16396 14424 16448
rect 15660 16396 15712 16448
rect 6103 16294 6155 16346
rect 6167 16294 6219 16346
rect 6231 16294 6283 16346
rect 6295 16294 6347 16346
rect 11224 16294 11276 16346
rect 11288 16294 11340 16346
rect 11352 16294 11404 16346
rect 11416 16294 11468 16346
rect 5356 16192 5408 16244
rect 5448 16235 5500 16244
rect 5448 16201 5457 16235
rect 5457 16201 5491 16235
rect 5491 16201 5500 16235
rect 5448 16192 5500 16201
rect 8116 16192 8168 16244
rect 9312 16192 9364 16244
rect 10416 16192 10468 16244
rect 15384 16235 15436 16244
rect 15384 16201 15393 16235
rect 15393 16201 15427 16235
rect 15427 16201 15436 16235
rect 15384 16192 15436 16201
rect 5632 16167 5684 16176
rect 3700 16099 3752 16108
rect 3700 16065 3709 16099
rect 3709 16065 3743 16099
rect 3743 16065 3752 16099
rect 3700 16056 3752 16065
rect 3976 16056 4028 16108
rect 5632 16133 5641 16167
rect 5641 16133 5675 16167
rect 5675 16133 5684 16167
rect 5632 16124 5684 16133
rect 4988 16056 5040 16108
rect 5816 16099 5868 16108
rect 5816 16065 5825 16099
rect 5825 16065 5859 16099
rect 5859 16065 5868 16099
rect 5816 16056 5868 16065
rect 6460 16056 6512 16108
rect 7104 16099 7156 16108
rect 7104 16065 7113 16099
rect 7113 16065 7147 16099
rect 7147 16065 7156 16099
rect 7104 16056 7156 16065
rect 8300 16124 8352 16176
rect 11060 16124 11112 16176
rect 8392 16056 8444 16108
rect 10324 16099 10376 16108
rect 7564 15988 7616 16040
rect 4068 15920 4120 15972
rect 7012 15963 7064 15972
rect 7012 15929 7021 15963
rect 7021 15929 7055 15963
rect 7055 15929 7064 15963
rect 7012 15920 7064 15929
rect 2504 15852 2556 15904
rect 3976 15895 4028 15904
rect 3976 15861 3985 15895
rect 3985 15861 4019 15895
rect 4019 15861 4028 15895
rect 3976 15852 4028 15861
rect 8208 15852 8260 15904
rect 10324 16065 10333 16099
rect 10333 16065 10367 16099
rect 10367 16065 10376 16099
rect 10324 16056 10376 16065
rect 11796 16099 11848 16108
rect 11796 16065 11805 16099
rect 11805 16065 11839 16099
rect 11839 16065 11848 16099
rect 11796 16056 11848 16065
rect 14372 16124 14424 16176
rect 15292 16167 15344 16176
rect 15292 16133 15301 16167
rect 15301 16133 15335 16167
rect 15335 16133 15344 16167
rect 15292 16124 15344 16133
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 12256 15988 12308 16040
rect 13176 16031 13228 16040
rect 13176 15997 13185 16031
rect 13185 15997 13219 16031
rect 13219 15997 13228 16031
rect 14464 16056 14516 16108
rect 15200 16099 15252 16108
rect 15200 16065 15209 16099
rect 15209 16065 15243 16099
rect 15243 16065 15252 16099
rect 15200 16056 15252 16065
rect 13176 15988 13228 15997
rect 15568 15988 15620 16040
rect 15660 16031 15712 16040
rect 15660 15997 15669 16031
rect 15669 15997 15703 16031
rect 15703 15997 15712 16031
rect 15660 15988 15712 15997
rect 10876 15920 10928 15972
rect 14740 15963 14792 15972
rect 14740 15929 14749 15963
rect 14749 15929 14783 15963
rect 14783 15929 14792 15963
rect 14740 15920 14792 15929
rect 3542 15750 3594 15802
rect 3606 15750 3658 15802
rect 3670 15750 3722 15802
rect 3734 15750 3786 15802
rect 8664 15750 8716 15802
rect 8728 15750 8780 15802
rect 8792 15750 8844 15802
rect 8856 15750 8908 15802
rect 13785 15750 13837 15802
rect 13849 15750 13901 15802
rect 13913 15750 13965 15802
rect 13977 15750 14029 15802
rect 1492 15648 1544 15700
rect 2504 15691 2556 15700
rect 2504 15657 2513 15691
rect 2513 15657 2547 15691
rect 2547 15657 2556 15691
rect 2504 15648 2556 15657
rect 10324 15648 10376 15700
rect 12992 15691 13044 15700
rect 2136 15580 2188 15632
rect 3332 15512 3384 15564
rect 2780 15444 2832 15496
rect 9220 15444 9272 15496
rect 10876 15487 10928 15496
rect 10876 15453 10885 15487
rect 10885 15453 10919 15487
rect 10919 15453 10928 15487
rect 10876 15444 10928 15453
rect 12532 15580 12584 15632
rect 12992 15657 13001 15691
rect 13001 15657 13035 15691
rect 13035 15657 13044 15691
rect 12992 15648 13044 15657
rect 13176 15691 13228 15700
rect 13176 15657 13185 15691
rect 13185 15657 13219 15691
rect 13219 15657 13228 15691
rect 13176 15648 13228 15657
rect 15200 15691 15252 15700
rect 15200 15657 15209 15691
rect 15209 15657 15243 15691
rect 15243 15657 15252 15691
rect 15200 15648 15252 15657
rect 15476 15580 15528 15632
rect 12256 15444 12308 15496
rect 14924 15487 14976 15496
rect 14924 15453 14933 15487
rect 14933 15453 14967 15487
rect 14967 15453 14976 15487
rect 14924 15444 14976 15453
rect 3148 15376 3200 15428
rect 4160 15419 4212 15428
rect 4160 15385 4169 15419
rect 4169 15385 4203 15419
rect 4203 15385 4212 15419
rect 4160 15376 4212 15385
rect 11060 15376 11112 15428
rect 12348 15376 12400 15428
rect 14096 15376 14148 15428
rect 2412 15308 2464 15360
rect 10324 15308 10376 15360
rect 14648 15308 14700 15360
rect 6103 15206 6155 15258
rect 6167 15206 6219 15258
rect 6231 15206 6283 15258
rect 6295 15206 6347 15258
rect 11224 15206 11276 15258
rect 11288 15206 11340 15258
rect 11352 15206 11404 15258
rect 11416 15206 11468 15258
rect 3976 15104 4028 15156
rect 6460 15147 6512 15156
rect 6460 15113 6469 15147
rect 6469 15113 6503 15147
rect 6503 15113 6512 15147
rect 6460 15104 6512 15113
rect 2412 15011 2464 15020
rect 2412 14977 2421 15011
rect 2421 14977 2455 15011
rect 2455 14977 2464 15011
rect 2412 14968 2464 14977
rect 3332 15011 3384 15020
rect 3332 14977 3341 15011
rect 3341 14977 3375 15011
rect 3375 14977 3384 15011
rect 3332 14968 3384 14977
rect 2136 14832 2188 14884
rect 4436 14943 4488 14952
rect 4436 14909 4445 14943
rect 4445 14909 4479 14943
rect 4479 14909 4488 14943
rect 4436 14900 4488 14909
rect 4988 14900 5040 14952
rect 7380 15036 7432 15088
rect 11888 15104 11940 15156
rect 12348 15104 12400 15156
rect 14924 15104 14976 15156
rect 11612 15036 11664 15088
rect 7564 14968 7616 15020
rect 11336 14968 11388 15020
rect 5448 14943 5500 14952
rect 5448 14909 5457 14943
rect 5457 14909 5491 14943
rect 5491 14909 5500 14943
rect 5448 14900 5500 14909
rect 4528 14832 4580 14884
rect 7288 14900 7340 14952
rect 8484 14943 8536 14952
rect 8484 14909 8493 14943
rect 8493 14909 8527 14943
rect 8527 14909 8536 14943
rect 11612 14943 11664 14952
rect 8484 14900 8536 14909
rect 11612 14909 11621 14943
rect 11621 14909 11655 14943
rect 11655 14909 11664 14943
rect 11612 14900 11664 14909
rect 12716 14968 12768 15020
rect 15016 15011 15068 15020
rect 11980 14943 12032 14952
rect 11980 14909 11989 14943
rect 11989 14909 12023 14943
rect 12023 14909 12032 14943
rect 11980 14900 12032 14909
rect 15016 14977 15025 15011
rect 15025 14977 15059 15011
rect 15059 14977 15068 15011
rect 15016 14968 15068 14977
rect 14004 14900 14056 14952
rect 14832 14900 14884 14952
rect 15016 14832 15068 14884
rect 2504 14764 2556 14816
rect 2964 14764 3016 14816
rect 12624 14764 12676 14816
rect 3542 14662 3594 14714
rect 3606 14662 3658 14714
rect 3670 14662 3722 14714
rect 3734 14662 3786 14714
rect 8664 14662 8716 14714
rect 8728 14662 8780 14714
rect 8792 14662 8844 14714
rect 8856 14662 8908 14714
rect 13785 14662 13837 14714
rect 13849 14662 13901 14714
rect 13913 14662 13965 14714
rect 13977 14662 14029 14714
rect 2780 14603 2832 14612
rect 2780 14569 2789 14603
rect 2789 14569 2823 14603
rect 2823 14569 2832 14603
rect 2780 14560 2832 14569
rect 4160 14560 4212 14612
rect 5448 14560 5500 14612
rect 7564 14603 7616 14612
rect 7564 14569 7573 14603
rect 7573 14569 7607 14603
rect 7607 14569 7616 14603
rect 7564 14560 7616 14569
rect 8484 14560 8536 14612
rect 11336 14603 11388 14612
rect 11336 14569 11345 14603
rect 11345 14569 11379 14603
rect 11379 14569 11388 14603
rect 11336 14560 11388 14569
rect 11980 14560 12032 14612
rect 14832 14603 14884 14612
rect 14832 14569 14841 14603
rect 14841 14569 14875 14603
rect 14875 14569 14884 14603
rect 14832 14560 14884 14569
rect 15292 14560 15344 14612
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 2964 14399 3016 14408
rect 2964 14365 2973 14399
rect 2973 14365 3007 14399
rect 3007 14365 3016 14399
rect 2964 14356 3016 14365
rect 3148 14399 3200 14408
rect 3148 14365 3157 14399
rect 3157 14365 3191 14399
rect 3191 14365 3200 14399
rect 3148 14356 3200 14365
rect 4160 14356 4212 14408
rect 4436 14399 4488 14408
rect 4436 14365 4445 14399
rect 4445 14365 4479 14399
rect 4479 14365 4488 14399
rect 4436 14356 4488 14365
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 4988 14356 5040 14408
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 8024 14356 8076 14408
rect 8300 14399 8352 14408
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 9220 14399 9272 14408
rect 9220 14365 9229 14399
rect 9229 14365 9263 14399
rect 9263 14365 9272 14399
rect 10968 14424 11020 14476
rect 9220 14356 9272 14365
rect 11612 14399 11664 14408
rect 11612 14365 11621 14399
rect 11621 14365 11655 14399
rect 11655 14365 11664 14399
rect 14188 14424 14240 14476
rect 11612 14356 11664 14365
rect 12440 14288 12492 14340
rect 1584 14220 1636 14272
rect 7196 14220 7248 14272
rect 10140 14220 10192 14272
rect 13268 14356 13320 14408
rect 14372 14288 14424 14340
rect 15660 14356 15712 14408
rect 15752 14331 15804 14340
rect 15752 14297 15761 14331
rect 15761 14297 15795 14331
rect 15795 14297 15804 14331
rect 15752 14288 15804 14297
rect 14556 14220 14608 14272
rect 6103 14118 6155 14170
rect 6167 14118 6219 14170
rect 6231 14118 6283 14170
rect 6295 14118 6347 14170
rect 11224 14118 11276 14170
rect 11288 14118 11340 14170
rect 11352 14118 11404 14170
rect 11416 14118 11468 14170
rect 2412 14016 2464 14068
rect 7288 14016 7340 14068
rect 8024 14059 8076 14068
rect 8024 14025 8033 14059
rect 8033 14025 8067 14059
rect 8067 14025 8076 14059
rect 8024 14016 8076 14025
rect 5540 13948 5592 14000
rect 1584 13923 1636 13932
rect 1584 13889 1593 13923
rect 1593 13889 1627 13923
rect 1627 13889 1636 13923
rect 1584 13880 1636 13889
rect 2964 13880 3016 13932
rect 3424 13880 3476 13932
rect 3792 13880 3844 13932
rect 3976 13880 4028 13932
rect 5080 13923 5132 13932
rect 5080 13889 5089 13923
rect 5089 13889 5123 13923
rect 5123 13889 5132 13923
rect 5080 13880 5132 13889
rect 5264 13880 5316 13932
rect 5356 13880 5408 13932
rect 7932 13923 7984 13932
rect 3240 13812 3292 13864
rect 7196 13855 7248 13864
rect 7196 13821 7205 13855
rect 7205 13821 7239 13855
rect 7239 13821 7248 13855
rect 7196 13812 7248 13821
rect 7932 13889 7941 13923
rect 7941 13889 7975 13923
rect 7975 13889 7984 13923
rect 7932 13880 7984 13889
rect 10968 14016 11020 14068
rect 11612 14016 11664 14068
rect 12900 14016 12952 14068
rect 13544 14016 13596 14068
rect 15568 14059 15620 14068
rect 15568 14025 15577 14059
rect 15577 14025 15611 14059
rect 15611 14025 15620 14059
rect 15568 14016 15620 14025
rect 11888 13991 11940 14000
rect 11888 13957 11897 13991
rect 11897 13957 11931 13991
rect 11931 13957 11940 13991
rect 11888 13948 11940 13957
rect 12440 13948 12492 14000
rect 13636 13948 13688 14000
rect 9588 13923 9640 13932
rect 9588 13889 9597 13923
rect 9597 13889 9631 13923
rect 9631 13889 9640 13923
rect 9588 13880 9640 13889
rect 11612 13880 11664 13932
rect 8300 13812 8352 13864
rect 9496 13855 9548 13864
rect 9496 13821 9505 13855
rect 9505 13821 9539 13855
rect 9539 13821 9548 13855
rect 9496 13812 9548 13821
rect 11152 13812 11204 13864
rect 11796 13923 11848 13932
rect 11796 13889 11805 13923
rect 11805 13889 11839 13923
rect 11839 13889 11848 13923
rect 11796 13880 11848 13889
rect 11980 13923 12032 13932
rect 11980 13889 12015 13923
rect 12015 13889 12032 13923
rect 11980 13880 12032 13889
rect 12900 13880 12952 13932
rect 14188 13923 14240 13932
rect 14188 13889 14197 13923
rect 14197 13889 14231 13923
rect 14231 13889 14240 13923
rect 14188 13880 14240 13889
rect 14372 13923 14424 13932
rect 14372 13889 14381 13923
rect 14381 13889 14415 13923
rect 14415 13889 14424 13923
rect 14372 13880 14424 13889
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 15660 13923 15712 13932
rect 15660 13889 15669 13923
rect 15669 13889 15703 13923
rect 15703 13889 15712 13923
rect 15660 13880 15712 13889
rect 15752 13923 15804 13932
rect 15752 13889 15761 13923
rect 15761 13889 15795 13923
rect 15795 13889 15804 13923
rect 15752 13880 15804 13889
rect 11612 13744 11664 13796
rect 14280 13812 14332 13864
rect 12348 13744 12400 13796
rect 2044 13719 2096 13728
rect 2044 13685 2053 13719
rect 2053 13685 2087 13719
rect 2087 13685 2096 13719
rect 2044 13676 2096 13685
rect 2596 13719 2648 13728
rect 2596 13685 2605 13719
rect 2605 13685 2639 13719
rect 2639 13685 2648 13719
rect 2596 13676 2648 13685
rect 4068 13676 4120 13728
rect 5172 13676 5224 13728
rect 9220 13676 9272 13728
rect 11336 13676 11388 13728
rect 11888 13676 11940 13728
rect 12072 13676 12124 13728
rect 12440 13676 12492 13728
rect 12716 13719 12768 13728
rect 12716 13685 12725 13719
rect 12725 13685 12759 13719
rect 12759 13685 12768 13719
rect 12716 13676 12768 13685
rect 3542 13574 3594 13626
rect 3606 13574 3658 13626
rect 3670 13574 3722 13626
rect 3734 13574 3786 13626
rect 8664 13574 8716 13626
rect 8728 13574 8780 13626
rect 8792 13574 8844 13626
rect 8856 13574 8908 13626
rect 13785 13574 13837 13626
rect 13849 13574 13901 13626
rect 13913 13574 13965 13626
rect 13977 13574 14029 13626
rect 2136 13515 2188 13524
rect 2136 13481 2145 13515
rect 2145 13481 2179 13515
rect 2179 13481 2188 13515
rect 2136 13472 2188 13481
rect 2596 13472 2648 13524
rect 3884 13472 3936 13524
rect 4988 13515 5040 13524
rect 4988 13481 4997 13515
rect 4997 13481 5031 13515
rect 5031 13481 5040 13515
rect 4988 13472 5040 13481
rect 8300 13472 8352 13524
rect 11060 13472 11112 13524
rect 12072 13472 12124 13524
rect 12348 13515 12400 13524
rect 12348 13481 12357 13515
rect 12357 13481 12391 13515
rect 12391 13481 12400 13515
rect 12348 13472 12400 13481
rect 14096 13472 14148 13524
rect 14188 13472 14240 13524
rect 9588 13404 9640 13456
rect 14832 13404 14884 13456
rect 11152 13379 11204 13388
rect 11152 13345 11161 13379
rect 11161 13345 11195 13379
rect 11195 13345 11204 13379
rect 11152 13336 11204 13345
rect 11796 13336 11848 13388
rect 2412 13268 2464 13320
rect 2872 13268 2924 13320
rect 3240 13311 3292 13320
rect 3240 13277 3249 13311
rect 3249 13277 3283 13311
rect 3283 13277 3292 13311
rect 3240 13268 3292 13277
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 4068 13311 4120 13320
rect 4068 13277 4077 13311
rect 4077 13277 4111 13311
rect 4111 13277 4120 13311
rect 4068 13268 4120 13277
rect 5080 13268 5132 13320
rect 5264 13311 5316 13320
rect 5264 13277 5273 13311
rect 5273 13277 5307 13311
rect 5307 13277 5316 13311
rect 5264 13268 5316 13277
rect 8760 13268 8812 13320
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9496 13311 9548 13320
rect 9220 13268 9272 13277
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 11336 13311 11388 13320
rect 5448 13200 5500 13252
rect 7840 13243 7892 13252
rect 7840 13209 7849 13243
rect 7849 13209 7883 13243
rect 7883 13209 7892 13243
rect 7840 13200 7892 13209
rect 9404 13200 9456 13252
rect 11336 13277 11345 13311
rect 11345 13277 11379 13311
rect 11379 13277 11388 13311
rect 11336 13268 11388 13277
rect 11060 13200 11112 13252
rect 12164 13243 12216 13252
rect 12164 13209 12173 13243
rect 12173 13209 12207 13243
rect 12207 13209 12216 13243
rect 12164 13200 12216 13209
rect 12440 13200 12492 13252
rect 13360 13243 13412 13252
rect 7196 13132 7248 13184
rect 8944 13175 8996 13184
rect 8944 13141 8953 13175
rect 8953 13141 8987 13175
rect 8987 13141 8996 13175
rect 8944 13132 8996 13141
rect 10692 13132 10744 13184
rect 13360 13209 13369 13243
rect 13369 13209 13403 13243
rect 13403 13209 13412 13243
rect 13360 13200 13412 13209
rect 13544 13200 13596 13252
rect 14280 13243 14332 13252
rect 14280 13209 14289 13243
rect 14289 13209 14323 13243
rect 14323 13209 14332 13243
rect 14280 13200 14332 13209
rect 14924 13243 14976 13252
rect 14924 13209 14933 13243
rect 14933 13209 14967 13243
rect 14967 13209 14976 13243
rect 14924 13200 14976 13209
rect 15108 13243 15160 13252
rect 15108 13209 15117 13243
rect 15117 13209 15151 13243
rect 15151 13209 15160 13243
rect 15108 13200 15160 13209
rect 15200 13132 15252 13184
rect 15476 13132 15528 13184
rect 6103 13030 6155 13082
rect 6167 13030 6219 13082
rect 6231 13030 6283 13082
rect 6295 13030 6347 13082
rect 11224 13030 11276 13082
rect 11288 13030 11340 13082
rect 11352 13030 11404 13082
rect 11416 13030 11468 13082
rect 3148 12928 3200 12980
rect 5264 12928 5316 12980
rect 5448 12928 5500 12980
rect 3056 12860 3108 12912
rect 4068 12903 4120 12912
rect 2044 12792 2096 12844
rect 1492 12724 1544 12776
rect 3424 12792 3476 12844
rect 4068 12869 4077 12903
rect 4077 12869 4111 12903
rect 4111 12869 4120 12903
rect 4068 12860 4120 12869
rect 3884 12792 3936 12844
rect 5264 12792 5316 12844
rect 8944 12928 8996 12980
rect 9128 12928 9180 12980
rect 7196 12903 7248 12912
rect 7196 12869 7205 12903
rect 7205 12869 7239 12903
rect 7239 12869 7248 12903
rect 7196 12860 7248 12869
rect 9312 12860 9364 12912
rect 10876 12928 10928 12980
rect 11980 12928 12032 12980
rect 12992 12928 13044 12980
rect 14372 12971 14424 12980
rect 14372 12937 14381 12971
rect 14381 12937 14415 12971
rect 14415 12937 14424 12971
rect 14372 12928 14424 12937
rect 15016 12971 15068 12980
rect 15016 12937 15025 12971
rect 15025 12937 15059 12971
rect 15059 12937 15068 12971
rect 15016 12928 15068 12937
rect 10692 12903 10744 12912
rect 10692 12869 10701 12903
rect 10701 12869 10735 12903
rect 10735 12869 10744 12903
rect 10692 12860 10744 12869
rect 11060 12860 11112 12912
rect 5172 12724 5224 12776
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 7656 12792 7708 12844
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 9680 12835 9732 12844
rect 9680 12801 9689 12835
rect 9689 12801 9723 12835
rect 9723 12801 9732 12835
rect 9680 12792 9732 12801
rect 11428 12792 11480 12844
rect 5356 12724 5408 12733
rect 8300 12767 8352 12776
rect 8300 12733 8309 12767
rect 8309 12733 8343 12767
rect 8343 12733 8352 12767
rect 8300 12724 8352 12733
rect 9864 12724 9916 12776
rect 12072 12792 12124 12844
rect 12440 12792 12492 12844
rect 12900 12835 12952 12844
rect 12900 12801 12909 12835
rect 12909 12801 12943 12835
rect 12943 12801 12952 12835
rect 12900 12792 12952 12801
rect 13360 12792 13412 12844
rect 14188 12835 14240 12844
rect 14188 12801 14197 12835
rect 14197 12801 14231 12835
rect 14231 12801 14240 12835
rect 14188 12792 14240 12801
rect 14372 12792 14424 12844
rect 15108 12792 15160 12844
rect 15476 12835 15528 12844
rect 15476 12801 15485 12835
rect 15485 12801 15519 12835
rect 15519 12801 15528 12835
rect 15476 12792 15528 12801
rect 15568 12792 15620 12844
rect 12624 12656 12676 12708
rect 13176 12656 13228 12708
rect 1860 12631 1912 12640
rect 1860 12597 1869 12631
rect 1869 12597 1903 12631
rect 1903 12597 1912 12631
rect 1860 12588 1912 12597
rect 2044 12588 2096 12640
rect 7472 12588 7524 12640
rect 9312 12588 9364 12640
rect 9496 12588 9548 12640
rect 15016 12588 15068 12640
rect 3542 12486 3594 12538
rect 3606 12486 3658 12538
rect 3670 12486 3722 12538
rect 3734 12486 3786 12538
rect 8664 12486 8716 12538
rect 8728 12486 8780 12538
rect 8792 12486 8844 12538
rect 8856 12486 8908 12538
rect 13785 12486 13837 12538
rect 13849 12486 13901 12538
rect 13913 12486 13965 12538
rect 13977 12486 14029 12538
rect 1676 12384 1728 12436
rect 1768 12316 1820 12368
rect 1952 12384 2004 12436
rect 4068 12384 4120 12436
rect 7288 12384 7340 12436
rect 7840 12384 7892 12436
rect 11428 12384 11480 12436
rect 12256 12427 12308 12436
rect 12256 12393 12265 12427
rect 12265 12393 12299 12427
rect 12299 12393 12308 12427
rect 12256 12384 12308 12393
rect 12716 12427 12768 12436
rect 12716 12393 12725 12427
rect 12725 12393 12759 12427
rect 12759 12393 12768 12427
rect 12716 12384 12768 12393
rect 14188 12384 14240 12436
rect 10600 12316 10652 12368
rect 2136 12248 2188 12300
rect 7656 12291 7708 12300
rect 7656 12257 7665 12291
rect 7665 12257 7699 12291
rect 7699 12257 7708 12291
rect 7656 12248 7708 12257
rect 1492 12180 1544 12232
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 2228 12223 2280 12232
rect 2228 12189 2237 12223
rect 2237 12189 2271 12223
rect 2271 12189 2280 12223
rect 2228 12180 2280 12189
rect 7196 12180 7248 12232
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 8300 12248 8352 12300
rect 7472 12180 7524 12189
rect 9680 12223 9732 12232
rect 5540 12112 5592 12164
rect 6000 12112 6052 12164
rect 9680 12189 9689 12223
rect 9689 12189 9723 12223
rect 9723 12189 9732 12223
rect 9680 12180 9732 12189
rect 9864 12223 9916 12232
rect 9864 12189 9873 12223
rect 9873 12189 9907 12223
rect 9907 12189 9916 12223
rect 9864 12180 9916 12189
rect 11060 12180 11112 12232
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 11980 12248 12032 12300
rect 13360 12248 13412 12300
rect 14464 12316 14516 12368
rect 14924 12384 14976 12436
rect 15660 12384 15712 12436
rect 14188 12291 14240 12300
rect 14188 12257 14197 12291
rect 14197 12257 14231 12291
rect 14231 12257 14240 12291
rect 14188 12248 14240 12257
rect 14648 12248 14700 12300
rect 12072 12180 12124 12232
rect 12440 12223 12492 12232
rect 12440 12189 12449 12223
rect 12449 12189 12483 12223
rect 12483 12189 12492 12223
rect 13176 12223 13228 12232
rect 12440 12180 12492 12189
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 13728 12180 13780 12232
rect 14372 12223 14424 12232
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15476 12180 15528 12189
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 9772 12112 9824 12164
rect 11428 12112 11480 12164
rect 8024 12044 8076 12096
rect 8392 12087 8444 12096
rect 8392 12053 8401 12087
rect 8401 12053 8435 12087
rect 8435 12053 8444 12087
rect 8392 12044 8444 12053
rect 14648 12044 14700 12096
rect 6103 11942 6155 11994
rect 6167 11942 6219 11994
rect 6231 11942 6283 11994
rect 6295 11942 6347 11994
rect 11224 11942 11276 11994
rect 11288 11942 11340 11994
rect 11352 11942 11404 11994
rect 11416 11942 11468 11994
rect 2872 11883 2924 11892
rect 2872 11849 2881 11883
rect 2881 11849 2915 11883
rect 2915 11849 2924 11883
rect 2872 11840 2924 11849
rect 3976 11883 4028 11892
rect 3976 11849 3985 11883
rect 3985 11849 4019 11883
rect 4019 11849 4028 11883
rect 3976 11840 4028 11849
rect 5172 11883 5224 11892
rect 5172 11849 5181 11883
rect 5181 11849 5215 11883
rect 5215 11849 5224 11883
rect 5172 11840 5224 11849
rect 7656 11840 7708 11892
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 9680 11840 9732 11849
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 13544 11840 13596 11892
rect 15752 11840 15804 11892
rect 2136 11772 2188 11824
rect 1768 11704 1820 11756
rect 2964 11636 3016 11688
rect 3424 11679 3476 11688
rect 2780 11568 2832 11620
rect 2872 11568 2924 11620
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 5632 11772 5684 11824
rect 6920 11704 6972 11756
rect 7932 11772 7984 11824
rect 7196 11704 7248 11756
rect 7472 11704 7524 11756
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 5724 11679 5776 11688
rect 4620 11636 4672 11645
rect 5724 11645 5733 11679
rect 5733 11645 5767 11679
rect 5767 11645 5776 11679
rect 5724 11636 5776 11645
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 8116 11568 8168 11620
rect 8392 11815 8444 11824
rect 8392 11781 8401 11815
rect 8401 11781 8435 11815
rect 8435 11781 8444 11815
rect 8392 11772 8444 11781
rect 9772 11772 9824 11824
rect 9496 11747 9548 11756
rect 9496 11713 9505 11747
rect 9505 11713 9539 11747
rect 9539 11713 9548 11747
rect 9496 11704 9548 11713
rect 14188 11772 14240 11824
rect 15108 11772 15160 11824
rect 10324 11704 10376 11756
rect 11612 11747 11664 11756
rect 11612 11713 11621 11747
rect 11621 11713 11655 11747
rect 11655 11713 11664 11747
rect 11612 11704 11664 11713
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 13084 11704 13136 11756
rect 13728 11747 13780 11756
rect 13728 11713 13737 11747
rect 13737 11713 13771 11747
rect 13771 11713 13780 11747
rect 13728 11704 13780 11713
rect 14004 11747 14056 11756
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 10692 11679 10744 11688
rect 10692 11645 10701 11679
rect 10701 11645 10735 11679
rect 10735 11645 10744 11679
rect 10692 11636 10744 11645
rect 11796 11636 11848 11688
rect 14924 11704 14976 11756
rect 8484 11568 8536 11620
rect 12072 11568 12124 11620
rect 13360 11568 13412 11620
rect 2136 11500 2188 11552
rect 8392 11500 8444 11552
rect 13636 11500 13688 11552
rect 14464 11636 14516 11688
rect 14924 11500 14976 11552
rect 15200 11543 15252 11552
rect 15200 11509 15209 11543
rect 15209 11509 15243 11543
rect 15243 11509 15252 11543
rect 15200 11500 15252 11509
rect 3542 11398 3594 11450
rect 3606 11398 3658 11450
rect 3670 11398 3722 11450
rect 3734 11398 3786 11450
rect 8664 11398 8716 11450
rect 8728 11398 8780 11450
rect 8792 11398 8844 11450
rect 8856 11398 8908 11450
rect 13785 11398 13837 11450
rect 13849 11398 13901 11450
rect 13913 11398 13965 11450
rect 13977 11398 14029 11450
rect 3424 11296 3476 11348
rect 1768 11160 1820 11212
rect 2136 11203 2188 11212
rect 2136 11169 2145 11203
rect 2145 11169 2179 11203
rect 2179 11169 2188 11203
rect 2136 11160 2188 11169
rect 1492 11092 1544 11144
rect 2044 11135 2096 11144
rect 2044 11101 2053 11135
rect 2053 11101 2087 11135
rect 2087 11101 2096 11135
rect 2872 11135 2924 11144
rect 2044 11092 2096 11101
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 5540 11228 5592 11280
rect 8392 11296 8444 11348
rect 9496 11296 9548 11348
rect 3884 11160 3936 11212
rect 4068 11135 4120 11144
rect 4068 11101 4077 11135
rect 4077 11101 4111 11135
rect 4111 11101 4120 11135
rect 4068 11092 4120 11101
rect 6920 11160 6972 11212
rect 8024 11228 8076 11280
rect 7380 11160 7432 11212
rect 10692 11160 10744 11212
rect 4620 11024 4672 11076
rect 2780 10956 2832 11008
rect 2872 10956 2924 11008
rect 6828 11024 6880 11076
rect 7104 11024 7156 11076
rect 7380 11067 7432 11076
rect 7380 11033 7415 11067
rect 7415 11033 7432 11067
rect 7380 11024 7432 11033
rect 7564 11024 7616 11076
rect 8484 11092 8536 11144
rect 9496 11092 9548 11144
rect 7656 10956 7708 11008
rect 8208 10956 8260 11008
rect 8392 10956 8444 11008
rect 9680 11024 9732 11076
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 10600 11135 10652 11144
rect 9864 11092 9916 11101
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 11980 11296 12032 11348
rect 12072 11296 12124 11348
rect 12992 11296 13044 11348
rect 13544 11296 13596 11348
rect 13636 11296 13688 11348
rect 11888 11228 11940 11280
rect 12808 11092 12860 11144
rect 14188 11160 14240 11212
rect 14096 11135 14148 11144
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 15476 11092 15528 11144
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 10048 10956 10100 11008
rect 10324 10956 10376 11008
rect 12440 11024 12492 11076
rect 12624 11024 12676 11076
rect 12532 10956 12584 11008
rect 13360 11024 13412 11076
rect 6103 10854 6155 10906
rect 6167 10854 6219 10906
rect 6231 10854 6283 10906
rect 6295 10854 6347 10906
rect 11224 10854 11276 10906
rect 11288 10854 11340 10906
rect 11352 10854 11404 10906
rect 11416 10854 11468 10906
rect 2780 10795 2832 10804
rect 2780 10761 2789 10795
rect 2789 10761 2823 10795
rect 2823 10761 2832 10795
rect 3884 10795 3936 10804
rect 2780 10752 2832 10761
rect 3884 10761 3893 10795
rect 3893 10761 3927 10795
rect 3927 10761 3936 10795
rect 3884 10752 3936 10761
rect 1952 10684 2004 10736
rect 2228 10659 2280 10668
rect 2228 10625 2237 10659
rect 2237 10625 2271 10659
rect 2271 10625 2280 10659
rect 2228 10616 2280 10625
rect 2412 10616 2464 10668
rect 4620 10752 4672 10804
rect 4528 10684 4580 10736
rect 7380 10752 7432 10804
rect 7472 10752 7524 10804
rect 8208 10752 8260 10804
rect 10416 10752 10468 10804
rect 10968 10795 11020 10804
rect 10968 10761 10977 10795
rect 10977 10761 11011 10795
rect 11011 10761 11020 10795
rect 10968 10752 11020 10761
rect 9404 10684 9456 10736
rect 11888 10752 11940 10804
rect 14280 10752 14332 10804
rect 15476 10795 15528 10804
rect 15476 10761 15485 10795
rect 15485 10761 15519 10795
rect 15519 10761 15528 10795
rect 15476 10752 15528 10761
rect 11796 10684 11848 10736
rect 4896 10616 4948 10668
rect 3240 10548 3292 10600
rect 5448 10659 5500 10668
rect 5448 10625 5457 10659
rect 5457 10625 5491 10659
rect 5491 10625 5500 10659
rect 5448 10616 5500 10625
rect 7104 10616 7156 10668
rect 8392 10616 8444 10668
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 10048 10616 10100 10668
rect 5080 10591 5132 10600
rect 5080 10557 5089 10591
rect 5089 10557 5123 10591
rect 5123 10557 5132 10591
rect 5080 10548 5132 10557
rect 7380 10548 7432 10600
rect 7748 10591 7800 10600
rect 7748 10557 7757 10591
rect 7757 10557 7791 10591
rect 7791 10557 7800 10591
rect 7748 10548 7800 10557
rect 8116 10548 8168 10600
rect 9128 10548 9180 10600
rect 9956 10591 10008 10600
rect 9956 10557 9965 10591
rect 9965 10557 9999 10591
rect 9999 10557 10008 10591
rect 9956 10548 10008 10557
rect 5632 10480 5684 10532
rect 1860 10412 1912 10464
rect 7196 10455 7248 10464
rect 7196 10421 7205 10455
rect 7205 10421 7239 10455
rect 7239 10421 7248 10455
rect 7196 10412 7248 10421
rect 7748 10412 7800 10464
rect 9036 10412 9088 10464
rect 10324 10480 10376 10532
rect 10876 10548 10928 10600
rect 11060 10616 11112 10668
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 12440 10616 12492 10668
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 12808 10548 12860 10600
rect 14372 10616 14424 10668
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 15108 10616 15160 10668
rect 13544 10480 13596 10532
rect 15200 10480 15252 10532
rect 10140 10412 10192 10464
rect 11796 10412 11848 10464
rect 3542 10310 3594 10362
rect 3606 10310 3658 10362
rect 3670 10310 3722 10362
rect 3734 10310 3786 10362
rect 8664 10310 8716 10362
rect 8728 10310 8780 10362
rect 8792 10310 8844 10362
rect 8856 10310 8908 10362
rect 13785 10310 13837 10362
rect 13849 10310 13901 10362
rect 13913 10310 13965 10362
rect 13977 10310 14029 10362
rect 2228 10208 2280 10260
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 7104 10208 7156 10260
rect 9772 10251 9824 10260
rect 9772 10217 9781 10251
rect 9781 10217 9815 10251
rect 9815 10217 9824 10251
rect 9772 10208 9824 10217
rect 9956 10208 10008 10260
rect 10784 10208 10836 10260
rect 10876 10208 10928 10260
rect 1952 10115 2004 10124
rect 1952 10081 1961 10115
rect 1961 10081 1995 10115
rect 1995 10081 2004 10115
rect 1952 10072 2004 10081
rect 2412 10072 2464 10124
rect 2872 10140 2924 10192
rect 6828 10140 6880 10192
rect 5908 10115 5960 10124
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 3056 10004 3108 10056
rect 3240 10047 3292 10056
rect 3240 10013 3249 10047
rect 3249 10013 3283 10047
rect 3283 10013 3292 10047
rect 3240 10004 3292 10013
rect 5908 10081 5917 10115
rect 5917 10081 5951 10115
rect 5951 10081 5960 10115
rect 5908 10072 5960 10081
rect 8024 10115 8076 10124
rect 8024 10081 8033 10115
rect 8033 10081 8067 10115
rect 8067 10081 8076 10115
rect 8024 10072 8076 10081
rect 9680 10140 9732 10192
rect 11980 10208 12032 10260
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 7932 10047 7984 10056
rect 5816 9936 5868 9988
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 8392 10047 8444 10056
rect 7472 9936 7524 9988
rect 7748 9936 7800 9988
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 9036 10004 9088 10056
rect 10324 10115 10376 10124
rect 10324 10081 10333 10115
rect 10333 10081 10367 10115
rect 10367 10081 10376 10115
rect 10324 10072 10376 10081
rect 10784 10072 10836 10124
rect 9864 9936 9916 9988
rect 2044 9868 2096 9920
rect 3240 9868 3292 9920
rect 7564 9868 7616 9920
rect 9128 9911 9180 9920
rect 9128 9877 9137 9911
rect 9137 9877 9171 9911
rect 9171 9877 9180 9911
rect 9128 9868 9180 9877
rect 9680 9868 9732 9920
rect 10140 9868 10192 9920
rect 11060 9936 11112 9988
rect 13084 10140 13136 10192
rect 14924 10072 14976 10124
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 14096 10047 14148 10056
rect 14096 10013 14105 10047
rect 14105 10013 14139 10047
rect 14139 10013 14148 10047
rect 14096 10004 14148 10013
rect 15108 10047 15160 10056
rect 15108 10013 15117 10047
rect 15117 10013 15151 10047
rect 15151 10013 15160 10047
rect 15108 10004 15160 10013
rect 11980 9979 12032 9988
rect 11980 9945 11989 9979
rect 11989 9945 12023 9979
rect 12023 9945 12032 9979
rect 11980 9936 12032 9945
rect 12440 9936 12492 9988
rect 12624 9936 12676 9988
rect 14188 9936 14240 9988
rect 14648 9936 14700 9988
rect 12992 9911 13044 9920
rect 12992 9877 13001 9911
rect 13001 9877 13035 9911
rect 13035 9877 13044 9911
rect 14464 9911 14516 9920
rect 12992 9868 13044 9877
rect 14464 9877 14473 9911
rect 14473 9877 14507 9911
rect 14507 9877 14516 9911
rect 14464 9868 14516 9877
rect 6103 9766 6155 9818
rect 6167 9766 6219 9818
rect 6231 9766 6283 9818
rect 6295 9766 6347 9818
rect 11224 9766 11276 9818
rect 11288 9766 11340 9818
rect 11352 9766 11404 9818
rect 11416 9766 11468 9818
rect 1952 9664 2004 9716
rect 7012 9664 7064 9716
rect 8116 9664 8168 9716
rect 9496 9664 9548 9716
rect 9772 9664 9824 9716
rect 2136 9571 2188 9580
rect 2136 9537 2144 9571
rect 2144 9537 2178 9571
rect 2178 9537 2188 9571
rect 2136 9528 2188 9537
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 3240 9528 3292 9580
rect 5908 9596 5960 9648
rect 9956 9664 10008 9716
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 5816 9503 5868 9512
rect 5816 9469 5825 9503
rect 5825 9469 5859 9503
rect 5859 9469 5868 9503
rect 5816 9460 5868 9469
rect 8392 9460 8444 9512
rect 9588 9528 9640 9580
rect 9956 9571 10008 9604
rect 9956 9552 9965 9571
rect 9965 9552 9999 9571
rect 9999 9552 10008 9571
rect 11704 9596 11756 9648
rect 14740 9596 14792 9648
rect 10600 9528 10652 9580
rect 11612 9528 11664 9580
rect 12532 9528 12584 9580
rect 12900 9528 12952 9580
rect 13544 9528 13596 9580
rect 14832 9571 14884 9580
rect 14832 9537 14841 9571
rect 14841 9537 14875 9571
rect 14875 9537 14884 9571
rect 14832 9528 14884 9537
rect 15200 9528 15252 9580
rect 15292 9571 15344 9580
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 2964 9392 3016 9444
rect 7196 9392 7248 9444
rect 8300 9392 8352 9444
rect 13084 9392 13136 9444
rect 13452 9392 13504 9444
rect 5724 9324 5776 9376
rect 6000 9324 6052 9376
rect 9680 9324 9732 9376
rect 10508 9324 10560 9376
rect 12716 9324 12768 9376
rect 14464 9460 14516 9512
rect 14740 9460 14792 9512
rect 14464 9324 14516 9376
rect 3542 9222 3594 9274
rect 3606 9222 3658 9274
rect 3670 9222 3722 9274
rect 3734 9222 3786 9274
rect 8664 9222 8716 9274
rect 8728 9222 8780 9274
rect 8792 9222 8844 9274
rect 8856 9222 8908 9274
rect 13785 9222 13837 9274
rect 13849 9222 13901 9274
rect 13913 9222 13965 9274
rect 13977 9222 14029 9274
rect 2136 9163 2188 9172
rect 2136 9129 2145 9163
rect 2145 9129 2179 9163
rect 2179 9129 2188 9163
rect 2136 9120 2188 9129
rect 4068 9120 4120 9172
rect 10232 9120 10284 9172
rect 11060 9120 11112 9172
rect 11612 9163 11664 9172
rect 11612 9129 11621 9163
rect 11621 9129 11655 9163
rect 11655 9129 11664 9163
rect 11612 9120 11664 9129
rect 13544 9163 13596 9172
rect 13544 9129 13553 9163
rect 13553 9129 13587 9163
rect 13587 9129 13596 9163
rect 13544 9120 13596 9129
rect 14556 9120 14608 9172
rect 5816 9052 5868 9104
rect 13452 9052 13504 9104
rect 4344 8984 4396 9036
rect 7564 8984 7616 9036
rect 7472 8959 7524 8968
rect 1860 8848 1912 8900
rect 1952 8891 2004 8900
rect 1952 8857 1961 8891
rect 1961 8857 1995 8891
rect 1995 8857 2004 8891
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 9128 8984 9180 9036
rect 10140 8984 10192 9036
rect 8300 8916 8352 8968
rect 9588 8916 9640 8968
rect 11980 8984 12032 9036
rect 12440 9027 12492 9036
rect 12440 8993 12449 9027
rect 12449 8993 12483 9027
rect 12483 8993 12492 9027
rect 12440 8984 12492 8993
rect 4436 8891 4488 8900
rect 1952 8848 2004 8857
rect 4436 8857 4445 8891
rect 4445 8857 4479 8891
rect 4479 8857 4488 8891
rect 4436 8848 4488 8857
rect 2872 8780 2924 8832
rect 7564 8891 7616 8900
rect 7564 8857 7573 8891
rect 7573 8857 7607 8891
rect 7607 8857 7616 8891
rect 7564 8848 7616 8857
rect 7748 8891 7800 8900
rect 7748 8857 7783 8891
rect 7783 8857 7800 8891
rect 7748 8848 7800 8857
rect 11520 8848 11572 8900
rect 14096 8916 14148 8968
rect 14740 8959 14792 8968
rect 12348 8848 12400 8900
rect 13452 8848 13504 8900
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 14924 8848 14976 8900
rect 15660 8891 15712 8900
rect 15660 8857 15669 8891
rect 15669 8857 15703 8891
rect 15703 8857 15712 8891
rect 15660 8848 15712 8857
rect 6103 8678 6155 8730
rect 6167 8678 6219 8730
rect 6231 8678 6283 8730
rect 6295 8678 6347 8730
rect 11224 8678 11276 8730
rect 11288 8678 11340 8730
rect 11352 8678 11404 8730
rect 11416 8678 11468 8730
rect 2228 8576 2280 8628
rect 3056 8576 3108 8628
rect 5080 8576 5132 8628
rect 7472 8576 7524 8628
rect 10324 8576 10376 8628
rect 13084 8619 13136 8628
rect 13084 8585 13093 8619
rect 13093 8585 13127 8619
rect 13127 8585 13136 8619
rect 13084 8576 13136 8585
rect 13176 8576 13228 8628
rect 13452 8619 13504 8628
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 2596 8483 2648 8492
rect 2596 8449 2605 8483
rect 2605 8449 2639 8483
rect 2639 8449 2648 8483
rect 6000 8508 6052 8560
rect 6920 8551 6972 8560
rect 6920 8517 6929 8551
rect 6929 8517 6963 8551
rect 6963 8517 6972 8551
rect 6920 8508 6972 8517
rect 2596 8440 2648 8449
rect 4620 8483 4672 8492
rect 1952 8372 2004 8424
rect 2412 8372 2464 8424
rect 2688 8372 2740 8424
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 4620 8440 4672 8449
rect 4436 8304 4488 8356
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 8116 8440 8168 8492
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 5816 8415 5868 8424
rect 5816 8381 5825 8415
rect 5825 8381 5859 8415
rect 5859 8381 5868 8415
rect 5816 8372 5868 8381
rect 7380 8372 7432 8424
rect 9036 8440 9088 8492
rect 11520 8508 11572 8560
rect 9956 8483 10008 8492
rect 9956 8449 9965 8483
rect 9965 8449 9999 8483
rect 9999 8449 10008 8483
rect 9956 8440 10008 8449
rect 8392 8415 8444 8424
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 8300 8347 8352 8356
rect 8300 8313 8309 8347
rect 8309 8313 8343 8347
rect 8343 8313 8352 8347
rect 8300 8304 8352 8313
rect 10508 8440 10560 8492
rect 12440 8508 12492 8560
rect 13636 8508 13688 8560
rect 12624 8440 12676 8492
rect 12900 8440 12952 8492
rect 14280 8483 14332 8492
rect 14280 8449 14289 8483
rect 14289 8449 14323 8483
rect 14323 8449 14332 8483
rect 14280 8440 14332 8449
rect 15200 8483 15252 8492
rect 15200 8449 15209 8483
rect 15209 8449 15243 8483
rect 15243 8449 15252 8483
rect 15200 8440 15252 8449
rect 12072 8415 12124 8424
rect 12072 8381 12081 8415
rect 12081 8381 12115 8415
rect 12115 8381 12124 8415
rect 12072 8372 12124 8381
rect 13268 8372 13320 8424
rect 6460 8236 6512 8288
rect 10876 8236 10928 8288
rect 12992 8304 13044 8356
rect 13360 8304 13412 8356
rect 15292 8372 15344 8424
rect 12716 8236 12768 8288
rect 13452 8236 13504 8288
rect 3542 8134 3594 8186
rect 3606 8134 3658 8186
rect 3670 8134 3722 8186
rect 3734 8134 3786 8186
rect 8664 8134 8716 8186
rect 8728 8134 8780 8186
rect 8792 8134 8844 8186
rect 8856 8134 8908 8186
rect 13785 8134 13837 8186
rect 13849 8134 13901 8186
rect 13913 8134 13965 8186
rect 13977 8134 14029 8186
rect 2596 8032 2648 8084
rect 6552 8032 6604 8084
rect 7380 8032 7432 8084
rect 8392 8032 8444 8084
rect 9680 8032 9732 8084
rect 10140 8032 10192 8084
rect 12348 8075 12400 8084
rect 8208 7964 8260 8016
rect 4620 7939 4672 7948
rect 4620 7905 4629 7939
rect 4629 7905 4663 7939
rect 4663 7905 4672 7939
rect 4620 7896 4672 7905
rect 2872 7828 2924 7880
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 5356 7871 5408 7880
rect 4712 7828 4764 7837
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 7380 7896 7432 7948
rect 6644 7871 6696 7880
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 7288 7828 7340 7880
rect 8116 7828 8168 7880
rect 9036 7964 9088 8016
rect 10692 7939 10744 7948
rect 10692 7905 10701 7939
rect 10701 7905 10735 7939
rect 10735 7905 10744 7939
rect 10692 7896 10744 7905
rect 12348 8041 12357 8075
rect 12357 8041 12391 8075
rect 12391 8041 12400 8075
rect 12348 8032 12400 8041
rect 14096 8075 14148 8084
rect 14096 8041 14105 8075
rect 14105 8041 14139 8075
rect 14139 8041 14148 8075
rect 14096 8032 14148 8041
rect 13636 7964 13688 8016
rect 15200 8032 15252 8084
rect 13360 7896 13412 7948
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 10048 7828 10100 7880
rect 10140 7828 10192 7880
rect 10876 7871 10928 7880
rect 10876 7837 10885 7871
rect 10885 7837 10919 7871
rect 10919 7837 10928 7871
rect 10876 7828 10928 7837
rect 13084 7828 13136 7880
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 15108 7964 15160 8016
rect 14372 7871 14424 7880
rect 14372 7837 14381 7871
rect 14381 7837 14415 7871
rect 14415 7837 14424 7871
rect 14648 7871 14700 7880
rect 14372 7828 14424 7837
rect 14648 7837 14657 7871
rect 14657 7837 14691 7871
rect 14691 7837 14700 7871
rect 14648 7828 14700 7837
rect 2780 7692 2832 7744
rect 5816 7760 5868 7812
rect 6736 7692 6788 7744
rect 7104 7692 7156 7744
rect 7564 7760 7616 7812
rect 8208 7760 8260 7812
rect 9404 7760 9456 7812
rect 11612 7803 11664 7812
rect 11612 7769 11621 7803
rect 11621 7769 11655 7803
rect 11655 7769 11664 7803
rect 11612 7760 11664 7769
rect 11888 7760 11940 7812
rect 12900 7760 12952 7812
rect 14832 7760 14884 7812
rect 15292 7803 15344 7812
rect 15292 7769 15301 7803
rect 15301 7769 15335 7803
rect 15335 7769 15344 7803
rect 15292 7760 15344 7769
rect 10600 7692 10652 7744
rect 12440 7692 12492 7744
rect 13084 7692 13136 7744
rect 13452 7692 13504 7744
rect 6103 7590 6155 7642
rect 6167 7590 6219 7642
rect 6231 7590 6283 7642
rect 6295 7590 6347 7642
rect 11224 7590 11276 7642
rect 11288 7590 11340 7642
rect 11352 7590 11404 7642
rect 11416 7590 11468 7642
rect 1860 7488 1912 7540
rect 2688 7420 2740 7472
rect 4620 7488 4672 7540
rect 6920 7488 6972 7540
rect 7472 7488 7524 7540
rect 2596 7352 2648 7404
rect 2780 7395 2832 7404
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 3976 7395 4028 7404
rect 2780 7352 2832 7361
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 7748 7463 7800 7472
rect 7748 7429 7757 7463
rect 7757 7429 7791 7463
rect 7791 7429 7800 7463
rect 7748 7420 7800 7429
rect 8392 7488 8444 7540
rect 9680 7488 9732 7540
rect 10140 7488 10192 7540
rect 2872 7284 2924 7336
rect 4804 7259 4856 7268
rect 4804 7225 4813 7259
rect 4813 7225 4847 7259
rect 4847 7225 4856 7259
rect 4804 7216 4856 7225
rect 5724 7284 5776 7336
rect 6736 7352 6788 7404
rect 7472 7352 7524 7404
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 7932 7352 7984 7404
rect 8484 7352 8536 7404
rect 10600 7420 10652 7472
rect 10048 7395 10100 7404
rect 10048 7361 10057 7395
rect 10057 7361 10091 7395
rect 10091 7361 10100 7395
rect 10048 7352 10100 7361
rect 10876 7395 10928 7404
rect 10876 7361 10885 7395
rect 10885 7361 10919 7395
rect 10919 7361 10928 7395
rect 10876 7352 10928 7361
rect 10968 7352 11020 7404
rect 12164 7488 12216 7540
rect 13820 7488 13872 7540
rect 14096 7488 14148 7540
rect 14740 7488 14792 7540
rect 15292 7488 15344 7540
rect 13176 7420 13228 7472
rect 5816 7216 5868 7268
rect 7012 7284 7064 7336
rect 7104 7216 7156 7268
rect 7472 7191 7524 7200
rect 7472 7157 7481 7191
rect 7481 7157 7515 7191
rect 7515 7157 7524 7191
rect 7472 7148 7524 7157
rect 8300 7284 8352 7336
rect 11060 7284 11112 7336
rect 11980 7352 12032 7404
rect 12072 7395 12124 7404
rect 12072 7361 12081 7395
rect 12081 7361 12115 7395
rect 12115 7361 12124 7395
rect 12072 7352 12124 7361
rect 12256 7352 12308 7404
rect 12716 7395 12768 7404
rect 12716 7361 12725 7395
rect 12725 7361 12759 7395
rect 12759 7361 12768 7395
rect 12716 7352 12768 7361
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 14740 7352 14792 7404
rect 15108 7352 15160 7404
rect 9036 7216 9088 7268
rect 12624 7284 12676 7336
rect 14372 7284 14424 7336
rect 8116 7148 8168 7200
rect 11612 7148 11664 7200
rect 11704 7148 11756 7200
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13360 7148 13412 7200
rect 14556 7148 14608 7200
rect 3542 7046 3594 7098
rect 3606 7046 3658 7098
rect 3670 7046 3722 7098
rect 3734 7046 3786 7098
rect 8664 7046 8716 7098
rect 8728 7046 8780 7098
rect 8792 7046 8844 7098
rect 8856 7046 8908 7098
rect 13785 7046 13837 7098
rect 13849 7046 13901 7098
rect 13913 7046 13965 7098
rect 13977 7046 14029 7098
rect 2412 6987 2464 6996
rect 2412 6953 2421 6987
rect 2421 6953 2455 6987
rect 2455 6953 2464 6987
rect 2412 6944 2464 6953
rect 2780 6944 2832 6996
rect 7472 6944 7524 6996
rect 7564 6944 7616 6996
rect 8024 6919 8076 6928
rect 3240 6740 3292 6792
rect 2872 6672 2924 6724
rect 3056 6715 3108 6724
rect 3056 6681 3065 6715
rect 3065 6681 3099 6715
rect 3099 6681 3108 6715
rect 4528 6808 4580 6860
rect 7104 6851 7156 6860
rect 7104 6817 7113 6851
rect 7113 6817 7147 6851
rect 7147 6817 7156 6851
rect 7104 6808 7156 6817
rect 4896 6740 4948 6792
rect 5448 6740 5500 6792
rect 5908 6740 5960 6792
rect 6644 6740 6696 6792
rect 6828 6783 6880 6792
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 8024 6885 8033 6919
rect 8033 6885 8067 6919
rect 8067 6885 8076 6919
rect 8024 6876 8076 6885
rect 3056 6672 3108 6681
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 1676 6604 1728 6656
rect 5356 6604 5408 6656
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 7472 6740 7524 6792
rect 8760 6808 8812 6860
rect 9404 6808 9456 6860
rect 7288 6604 7340 6656
rect 7656 6604 7708 6656
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 10692 6876 10744 6928
rect 11060 6944 11112 6996
rect 12072 6944 12124 6996
rect 13176 6876 13228 6928
rect 10324 6808 10376 6860
rect 10876 6672 10928 6724
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 13544 6808 13596 6860
rect 11796 6740 11848 6749
rect 14372 6808 14424 6860
rect 15384 6808 15436 6860
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 11428 6672 11480 6724
rect 13176 6672 13228 6724
rect 14280 6672 14332 6724
rect 8024 6604 8076 6656
rect 10968 6604 11020 6656
rect 11796 6604 11848 6656
rect 13084 6604 13136 6656
rect 15016 6647 15068 6656
rect 15016 6613 15025 6647
rect 15025 6613 15059 6647
rect 15059 6613 15068 6647
rect 15016 6604 15068 6613
rect 6103 6502 6155 6554
rect 6167 6502 6219 6554
rect 6231 6502 6283 6554
rect 6295 6502 6347 6554
rect 11224 6502 11276 6554
rect 11288 6502 11340 6554
rect 11352 6502 11404 6554
rect 11416 6502 11468 6554
rect 3240 6443 3292 6452
rect 3240 6409 3249 6443
rect 3249 6409 3283 6443
rect 3283 6409 3292 6443
rect 3240 6400 3292 6409
rect 4896 6443 4948 6452
rect 1584 6332 1636 6384
rect 4896 6409 4905 6443
rect 4905 6409 4939 6443
rect 4939 6409 4948 6443
rect 4896 6400 4948 6409
rect 5448 6400 5500 6452
rect 7932 6400 7984 6452
rect 8208 6400 8260 6452
rect 8760 6443 8812 6452
rect 8760 6409 8769 6443
rect 8769 6409 8803 6443
rect 8803 6409 8812 6443
rect 8760 6400 8812 6409
rect 12072 6443 12124 6452
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 3792 6239 3844 6248
rect 3792 6205 3801 6239
rect 3801 6205 3835 6239
rect 3835 6205 3844 6239
rect 3792 6196 3844 6205
rect 9680 6332 9732 6384
rect 6552 6307 6604 6316
rect 4436 6196 4488 6248
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 6828 6264 6880 6316
rect 5448 6239 5500 6248
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 5448 6196 5500 6205
rect 5540 6239 5592 6248
rect 5540 6205 5549 6239
rect 5549 6205 5583 6239
rect 5583 6205 5592 6239
rect 5540 6196 5592 6205
rect 6644 6196 6696 6248
rect 7012 6239 7064 6248
rect 7012 6205 7021 6239
rect 7021 6205 7055 6239
rect 7055 6205 7064 6239
rect 7012 6196 7064 6205
rect 7840 6264 7892 6316
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 8392 6264 8444 6316
rect 8300 6196 8352 6248
rect 8484 6196 8536 6248
rect 9772 6264 9824 6316
rect 10692 6332 10744 6384
rect 11428 6332 11480 6384
rect 10784 6264 10836 6316
rect 12072 6409 12081 6443
rect 12081 6409 12115 6443
rect 12115 6409 12124 6443
rect 12072 6400 12124 6409
rect 12164 6400 12216 6452
rect 14648 6400 14700 6452
rect 12900 6332 12952 6384
rect 14464 6332 14516 6384
rect 12348 6264 12400 6316
rect 12808 6264 12860 6316
rect 13176 6264 13228 6316
rect 13544 6307 13596 6316
rect 13544 6273 13553 6307
rect 13553 6273 13587 6307
rect 13587 6273 13596 6307
rect 13544 6264 13596 6273
rect 13728 6264 13780 6316
rect 14924 6307 14976 6316
rect 14924 6273 14933 6307
rect 14933 6273 14967 6307
rect 14967 6273 14976 6307
rect 14924 6264 14976 6273
rect 15384 6307 15436 6316
rect 10324 6239 10376 6248
rect 10324 6205 10333 6239
rect 10333 6205 10367 6239
rect 10367 6205 10376 6239
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 10324 6196 10376 6205
rect 15292 6196 15344 6248
rect 2780 6128 2832 6180
rect 9772 6128 9824 6180
rect 14280 6171 14332 6180
rect 14280 6137 14289 6171
rect 14289 6137 14323 6171
rect 14323 6137 14332 6171
rect 14280 6128 14332 6137
rect 5448 6060 5500 6112
rect 3542 5958 3594 6010
rect 3606 5958 3658 6010
rect 3670 5958 3722 6010
rect 3734 5958 3786 6010
rect 8664 5958 8716 6010
rect 8728 5958 8780 6010
rect 8792 5958 8844 6010
rect 8856 5958 8908 6010
rect 13785 5958 13837 6010
rect 13849 5958 13901 6010
rect 13913 5958 13965 6010
rect 13977 5958 14029 6010
rect 3884 5856 3936 5908
rect 4436 5856 4488 5908
rect 5540 5856 5592 5908
rect 10784 5899 10836 5908
rect 10784 5865 10793 5899
rect 10793 5865 10827 5899
rect 10827 5865 10836 5899
rect 10784 5856 10836 5865
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 1860 5652 1912 5704
rect 2780 5652 2832 5704
rect 3056 5788 3108 5840
rect 3240 5788 3292 5840
rect 5448 5788 5500 5840
rect 7012 5788 7064 5840
rect 7656 5788 7708 5840
rect 4528 5695 4580 5704
rect 4528 5661 4537 5695
rect 4537 5661 4571 5695
rect 4571 5661 4580 5695
rect 4712 5695 4764 5704
rect 4528 5652 4580 5661
rect 4712 5661 4723 5695
rect 4723 5661 4764 5695
rect 4712 5652 4764 5661
rect 7932 5763 7984 5772
rect 7932 5729 7941 5763
rect 7941 5729 7975 5763
rect 7975 5729 7984 5763
rect 7932 5720 7984 5729
rect 8208 5788 8260 5840
rect 13360 5831 13412 5840
rect 13360 5797 13369 5831
rect 13369 5797 13403 5831
rect 13403 5797 13412 5831
rect 13360 5788 13412 5797
rect 14740 5788 14792 5840
rect 5080 5652 5132 5704
rect 5908 5652 5960 5704
rect 6736 5652 6788 5704
rect 7564 5652 7616 5704
rect 4068 5584 4120 5636
rect 6460 5584 6512 5636
rect 7472 5584 7524 5636
rect 1400 5516 1452 5568
rect 2136 5559 2188 5568
rect 2136 5525 2145 5559
rect 2145 5525 2179 5559
rect 2179 5525 2188 5559
rect 2136 5516 2188 5525
rect 3424 5516 3476 5568
rect 5724 5559 5776 5568
rect 5724 5525 5733 5559
rect 5733 5525 5767 5559
rect 5767 5525 5776 5559
rect 5724 5516 5776 5525
rect 6552 5516 6604 5568
rect 8300 5652 8352 5704
rect 8392 5652 8444 5704
rect 8484 5584 8536 5636
rect 9864 5652 9916 5704
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 10968 5584 11020 5636
rect 13452 5652 13504 5704
rect 13728 5652 13780 5704
rect 12440 5584 12492 5636
rect 13544 5584 13596 5636
rect 8208 5516 8260 5568
rect 10416 5559 10468 5568
rect 10416 5525 10425 5559
rect 10425 5525 10459 5559
rect 10459 5525 10468 5559
rect 10416 5516 10468 5525
rect 10508 5516 10560 5568
rect 10692 5516 10744 5568
rect 12164 5516 12216 5568
rect 12348 5516 12400 5568
rect 12992 5559 13044 5568
rect 12992 5525 13001 5559
rect 13001 5525 13035 5559
rect 13035 5525 13044 5559
rect 12992 5516 13044 5525
rect 14832 5720 14884 5772
rect 15016 5763 15068 5772
rect 15016 5729 15025 5763
rect 15025 5729 15059 5763
rect 15059 5729 15068 5763
rect 15016 5720 15068 5729
rect 14372 5652 14424 5704
rect 14556 5652 14608 5704
rect 15108 5652 15160 5704
rect 14648 5584 14700 5636
rect 15384 5584 15436 5636
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 15200 5516 15252 5568
rect 6103 5414 6155 5466
rect 6167 5414 6219 5466
rect 6231 5414 6283 5466
rect 6295 5414 6347 5466
rect 11224 5414 11276 5466
rect 11288 5414 11340 5466
rect 11352 5414 11404 5466
rect 11416 5414 11468 5466
rect 2780 5312 2832 5364
rect 3332 5312 3384 5364
rect 6736 5312 6788 5364
rect 7564 5312 7616 5364
rect 8208 5312 8260 5364
rect 10416 5355 10468 5364
rect 10416 5321 10425 5355
rect 10425 5321 10459 5355
rect 10459 5321 10468 5355
rect 10416 5312 10468 5321
rect 10508 5355 10560 5364
rect 10508 5321 10517 5355
rect 10517 5321 10551 5355
rect 10551 5321 10560 5355
rect 10508 5312 10560 5321
rect 3976 5244 4028 5296
rect 1768 5176 1820 5228
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 3424 5219 3476 5228
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 5080 5244 5132 5296
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 5540 5219 5592 5228
rect 4988 5083 5040 5092
rect 4988 5049 4997 5083
rect 4997 5049 5031 5083
rect 5031 5049 5040 5083
rect 4988 5040 5040 5049
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 5632 5176 5684 5228
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 7012 5176 7064 5228
rect 7472 5176 7524 5228
rect 7840 5219 7892 5228
rect 7840 5185 7849 5219
rect 7849 5185 7883 5219
rect 7883 5185 7892 5219
rect 7840 5176 7892 5185
rect 9864 5244 9916 5296
rect 12440 5312 12492 5364
rect 12900 5355 12952 5364
rect 12900 5321 12909 5355
rect 12909 5321 12943 5355
rect 12943 5321 12952 5355
rect 12900 5312 12952 5321
rect 13544 5312 13596 5364
rect 14924 5312 14976 5364
rect 10600 5219 10652 5228
rect 10600 5185 10609 5219
rect 10609 5185 10643 5219
rect 10643 5185 10652 5219
rect 11796 5219 11848 5228
rect 10600 5176 10652 5185
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 11796 5176 11848 5185
rect 11980 5176 12032 5228
rect 12440 5176 12492 5228
rect 6644 5108 6696 5160
rect 7656 5108 7708 5160
rect 8300 5108 8352 5160
rect 10692 5108 10744 5160
rect 11612 5108 11664 5160
rect 11704 5108 11756 5160
rect 5356 5040 5408 5092
rect 6828 5040 6880 5092
rect 8208 5040 8260 5092
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 1676 4972 1728 5024
rect 2872 4972 2924 5024
rect 5080 4972 5132 5024
rect 8024 5015 8076 5024
rect 8024 4981 8033 5015
rect 8033 4981 8067 5015
rect 8067 4981 8076 5015
rect 8024 4972 8076 4981
rect 8300 4972 8352 5024
rect 10968 5040 11020 5092
rect 12256 5040 12308 5092
rect 10876 4972 10928 5024
rect 12900 5108 12952 5160
rect 13360 5151 13412 5160
rect 13360 5117 13369 5151
rect 13369 5117 13403 5151
rect 13403 5117 13412 5151
rect 13360 5108 13412 5117
rect 13912 5287 13964 5296
rect 13912 5253 13921 5287
rect 13921 5253 13955 5287
rect 13955 5253 13964 5287
rect 13912 5244 13964 5253
rect 13820 5176 13872 5228
rect 15108 5176 15160 5228
rect 14556 5108 14608 5160
rect 14188 4972 14240 5024
rect 3542 4870 3594 4922
rect 3606 4870 3658 4922
rect 3670 4870 3722 4922
rect 3734 4870 3786 4922
rect 8664 4870 8716 4922
rect 8728 4870 8780 4922
rect 8792 4870 8844 4922
rect 8856 4870 8908 4922
rect 13785 4870 13837 4922
rect 13849 4870 13901 4922
rect 13913 4870 13965 4922
rect 13977 4870 14029 4922
rect 1584 4768 1636 4820
rect 5172 4768 5224 4820
rect 7840 4768 7892 4820
rect 8392 4811 8444 4820
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 10140 4768 10192 4820
rect 11704 4811 11756 4820
rect 11704 4777 11713 4811
rect 11713 4777 11747 4811
rect 11747 4777 11756 4811
rect 11704 4768 11756 4777
rect 13176 4811 13228 4820
rect 13176 4777 13185 4811
rect 13185 4777 13219 4811
rect 13219 4777 13228 4811
rect 13176 4768 13228 4777
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 1768 4564 1820 4616
rect 1952 4607 2004 4616
rect 1952 4573 1961 4607
rect 1961 4573 1995 4607
rect 1995 4573 2004 4607
rect 1952 4564 2004 4573
rect 4804 4700 4856 4752
rect 5448 4700 5500 4752
rect 3424 4632 3476 4684
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5356 4607 5408 4616
rect 5080 4564 5132 4573
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 5908 4564 5960 4616
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 13268 4700 13320 4752
rect 13544 4700 13596 4752
rect 8300 4564 8352 4616
rect 8944 4607 8996 4616
rect 8944 4573 8953 4607
rect 8953 4573 8987 4607
rect 8987 4573 8996 4607
rect 8944 4564 8996 4573
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 10876 4564 10928 4616
rect 2320 4496 2372 4548
rect 2964 4428 3016 4480
rect 4068 4496 4120 4548
rect 5724 4496 5776 4548
rect 9312 4496 9364 4548
rect 10784 4539 10836 4548
rect 10784 4505 10793 4539
rect 10793 4505 10827 4539
rect 10827 4505 10836 4539
rect 10784 4496 10836 4505
rect 11060 4496 11112 4548
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 14188 4768 14240 4820
rect 15016 4632 15068 4684
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 14372 4564 14424 4616
rect 14648 4564 14700 4616
rect 11980 4496 12032 4548
rect 12716 4496 12768 4548
rect 12900 4496 12952 4548
rect 14740 4496 14792 4548
rect 5172 4428 5224 4480
rect 8116 4428 8168 4480
rect 8944 4428 8996 4480
rect 12440 4428 12492 4480
rect 15016 4428 15068 4480
rect 6103 4326 6155 4378
rect 6167 4326 6219 4378
rect 6231 4326 6283 4378
rect 6295 4326 6347 4378
rect 11224 4326 11276 4378
rect 11288 4326 11340 4378
rect 11352 4326 11404 4378
rect 11416 4326 11468 4378
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 2872 4131 2924 4140
rect 1584 4020 1636 4072
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 4528 4224 4580 4276
rect 4896 4267 4948 4276
rect 4896 4233 4905 4267
rect 4905 4233 4939 4267
rect 4939 4233 4948 4267
rect 4896 4224 4948 4233
rect 8024 4224 8076 4276
rect 5356 4088 5408 4140
rect 7840 4156 7892 4208
rect 4344 4020 4396 4072
rect 5448 4020 5500 4072
rect 6736 4088 6788 4140
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 7196 4088 7248 4140
rect 12440 4224 12492 4276
rect 15292 4224 15344 4276
rect 9220 4156 9272 4208
rect 6828 4020 6880 4072
rect 7748 4020 7800 4072
rect 9404 4088 9456 4140
rect 10784 4131 10836 4140
rect 10784 4097 10793 4131
rect 10793 4097 10827 4131
rect 10827 4097 10836 4131
rect 10784 4088 10836 4097
rect 12716 4156 12768 4208
rect 14372 4199 14424 4208
rect 14372 4165 14381 4199
rect 14381 4165 14415 4199
rect 14415 4165 14424 4199
rect 14372 4156 14424 4165
rect 14556 4199 14608 4208
rect 14556 4165 14565 4199
rect 14565 4165 14599 4199
rect 14599 4165 14608 4199
rect 14556 4156 14608 4165
rect 14924 4156 14976 4208
rect 15200 4199 15252 4208
rect 15200 4165 15209 4199
rect 15209 4165 15243 4199
rect 15243 4165 15252 4199
rect 15200 4156 15252 4165
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 12440 4088 12492 4140
rect 12532 4088 12584 4140
rect 12992 4088 13044 4140
rect 14280 4088 14332 4140
rect 6092 3952 6144 4004
rect 6920 3952 6972 4004
rect 8484 3952 8536 4004
rect 1768 3884 1820 3936
rect 4712 3884 4764 3936
rect 4804 3884 4856 3936
rect 8024 3884 8076 3936
rect 9496 4020 9548 4072
rect 12716 4020 12768 4072
rect 10784 3952 10836 4004
rect 14832 4020 14884 4072
rect 12900 3952 12952 4004
rect 13452 3952 13504 4004
rect 14464 3952 14516 4004
rect 9680 3884 9732 3936
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 11060 3884 11112 3936
rect 11152 3884 11204 3936
rect 12532 3884 12584 3936
rect 14188 3927 14240 3936
rect 14188 3893 14197 3927
rect 14197 3893 14231 3927
rect 14231 3893 14240 3927
rect 14188 3884 14240 3893
rect 3542 3782 3594 3834
rect 3606 3782 3658 3834
rect 3670 3782 3722 3834
rect 3734 3782 3786 3834
rect 8664 3782 8716 3834
rect 8728 3782 8780 3834
rect 8792 3782 8844 3834
rect 8856 3782 8908 3834
rect 13785 3782 13837 3834
rect 13849 3782 13901 3834
rect 13913 3782 13965 3834
rect 13977 3782 14029 3834
rect 1952 3544 2004 3596
rect 2320 3544 2372 3596
rect 4344 3612 4396 3664
rect 4528 3612 4580 3664
rect 5724 3612 5776 3664
rect 5908 3612 5960 3664
rect 7104 3680 7156 3732
rect 8300 3680 8352 3732
rect 9128 3680 9180 3732
rect 9496 3723 9548 3732
rect 9496 3689 9505 3723
rect 9505 3689 9539 3723
rect 9539 3689 9548 3723
rect 9496 3680 9548 3689
rect 12808 3680 12860 3732
rect 13544 3680 13596 3732
rect 14280 3680 14332 3732
rect 15384 3680 15436 3732
rect 8024 3612 8076 3664
rect 3148 3544 3200 3596
rect 8484 3612 8536 3664
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 1860 3476 1912 3528
rect 3884 3519 3936 3528
rect 3884 3485 3926 3519
rect 3926 3485 3936 3519
rect 3884 3476 3936 3485
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5908 3519 5960 3528
rect 5632 3476 5684 3485
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 6092 3476 6144 3528
rect 6736 3476 6788 3528
rect 5264 3408 5316 3460
rect 6828 3451 6880 3460
rect 3516 3340 3568 3392
rect 4068 3340 4120 3392
rect 5448 3340 5500 3392
rect 6828 3417 6837 3451
rect 6837 3417 6871 3451
rect 6871 3417 6880 3451
rect 6828 3408 6880 3417
rect 7196 3408 7248 3460
rect 9404 3544 9456 3596
rect 10324 3612 10376 3664
rect 11796 3612 11848 3664
rect 12624 3612 12676 3664
rect 8208 3476 8260 3528
rect 8668 3476 8720 3528
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 11152 3476 11204 3528
rect 11520 3544 11572 3596
rect 12164 3544 12216 3596
rect 12348 3476 12400 3528
rect 14188 3544 14240 3596
rect 12716 3408 12768 3460
rect 6000 3340 6052 3392
rect 6552 3340 6604 3392
rect 8392 3340 8444 3392
rect 9312 3340 9364 3392
rect 12808 3340 12860 3392
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14832 3544 14884 3596
rect 14280 3476 14332 3485
rect 15108 3476 15160 3528
rect 13820 3340 13872 3392
rect 13912 3340 13964 3392
rect 14464 3451 14516 3460
rect 14464 3417 14473 3451
rect 14473 3417 14507 3451
rect 14507 3417 14516 3451
rect 14464 3408 14516 3417
rect 14924 3340 14976 3392
rect 6103 3238 6155 3290
rect 6167 3238 6219 3290
rect 6231 3238 6283 3290
rect 6295 3238 6347 3290
rect 11224 3238 11276 3290
rect 11288 3238 11340 3290
rect 11352 3238 11404 3290
rect 11416 3238 11468 3290
rect 2596 3179 2648 3188
rect 2596 3145 2605 3179
rect 2605 3145 2639 3179
rect 2639 3145 2648 3179
rect 2596 3136 2648 3145
rect 4068 3136 4120 3188
rect 5264 3136 5316 3188
rect 1400 3111 1452 3120
rect 1400 3077 1409 3111
rect 1409 3077 1443 3111
rect 1443 3077 1452 3111
rect 3332 3111 3384 3120
rect 1400 3068 1452 3077
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 3332 3077 3341 3111
rect 3341 3077 3375 3111
rect 3375 3077 3384 3111
rect 3332 3068 3384 3077
rect 2688 3041 2740 3052
rect 2688 3007 2697 3041
rect 2697 3007 2731 3041
rect 2731 3007 2740 3041
rect 3148 3043 3200 3052
rect 2688 3000 2740 3007
rect 3148 3009 3157 3043
rect 3157 3009 3191 3043
rect 3191 3009 3200 3043
rect 3148 3000 3200 3009
rect 3516 3000 3568 3052
rect 7288 3068 7340 3120
rect 2136 2932 2188 2984
rect 5908 3000 5960 3052
rect 7840 3000 7892 3052
rect 9128 3136 9180 3188
rect 11520 3136 11572 3188
rect 8760 3068 8812 3120
rect 13176 3136 13228 3188
rect 17500 3136 17552 3188
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 8668 3043 8720 3052
rect 8668 3009 8677 3043
rect 8677 3009 8711 3043
rect 8711 3009 8720 3043
rect 9680 3043 9732 3052
rect 8668 3000 8720 3009
rect 9680 3009 9689 3043
rect 9689 3009 9723 3043
rect 9723 3009 9732 3043
rect 9680 3000 9732 3009
rect 12532 3068 12584 3120
rect 12808 3068 12860 3120
rect 13452 3068 13504 3120
rect 13544 3068 13596 3120
rect 13912 3111 13964 3120
rect 10508 3043 10560 3052
rect 10508 3009 10517 3043
rect 10517 3009 10551 3043
rect 10551 3009 10560 3043
rect 10508 3000 10560 3009
rect 11060 3000 11112 3052
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 13268 3000 13320 3052
rect 13912 3077 13921 3111
rect 13921 3077 13955 3111
rect 13955 3077 13964 3111
rect 13912 3068 13964 3077
rect 4436 2975 4488 2984
rect 4436 2941 4445 2975
rect 4445 2941 4479 2975
rect 4479 2941 4488 2975
rect 4436 2932 4488 2941
rect 4068 2864 4120 2916
rect 4252 2864 4304 2916
rect 5540 2932 5592 2984
rect 6000 2932 6052 2984
rect 6736 2932 6788 2984
rect 6828 2932 6880 2984
rect 7104 2975 7156 2984
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 9864 2975 9916 2984
rect 1860 2796 1912 2848
rect 3884 2796 3936 2848
rect 7012 2864 7064 2916
rect 9864 2941 9873 2975
rect 9873 2941 9907 2975
rect 9907 2941 9916 2975
rect 9864 2932 9916 2941
rect 9956 2932 10008 2984
rect 12900 2932 12952 2984
rect 13820 2932 13872 2984
rect 14096 3068 14148 3120
rect 14832 3111 14884 3120
rect 7748 2864 7800 2916
rect 7104 2796 7156 2848
rect 8392 2864 8444 2916
rect 9220 2864 9272 2916
rect 13176 2796 13228 2848
rect 13268 2796 13320 2848
rect 13452 2796 13504 2848
rect 14832 3077 14841 3111
rect 14841 3077 14875 3111
rect 14875 3077 14884 3111
rect 14832 3068 14884 3077
rect 15384 3000 15436 3052
rect 15752 2907 15804 2916
rect 15752 2873 15761 2907
rect 15761 2873 15795 2907
rect 15795 2873 15804 2907
rect 15752 2864 15804 2873
rect 3542 2694 3594 2746
rect 3606 2694 3658 2746
rect 3670 2694 3722 2746
rect 3734 2694 3786 2746
rect 8664 2694 8716 2746
rect 8728 2694 8780 2746
rect 8792 2694 8844 2746
rect 8856 2694 8908 2746
rect 13785 2694 13837 2746
rect 13849 2694 13901 2746
rect 13913 2694 13965 2746
rect 13977 2694 14029 2746
rect 5908 2592 5960 2644
rect 6920 2592 6972 2644
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 4712 2524 4764 2576
rect 8300 2592 8352 2644
rect 9864 2592 9916 2644
rect 2044 2456 2096 2508
rect 4804 2456 4856 2508
rect 20 2388 72 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2964 2388 3016 2440
rect 4068 2388 4120 2440
rect 5632 2456 5684 2508
rect 5448 2388 5500 2440
rect 5816 2388 5868 2440
rect 6552 2456 6604 2508
rect 8300 2456 8352 2508
rect 9404 2524 9456 2576
rect 11796 2592 11848 2644
rect 12716 2592 12768 2644
rect 14648 2592 14700 2644
rect 10048 2524 10100 2576
rect 1860 2320 1912 2372
rect 3884 2320 3936 2372
rect 5540 2320 5592 2372
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 7564 2431 7616 2440
rect 6736 2388 6788 2397
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 7564 2388 7616 2397
rect 8024 2431 8076 2440
rect 8024 2397 8033 2431
rect 8033 2397 8067 2431
rect 8067 2397 8076 2431
rect 8024 2388 8076 2397
rect 9128 2431 9180 2440
rect 7104 2320 7156 2372
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9956 2431 10008 2440
rect 9404 2320 9456 2372
rect 5632 2295 5684 2304
rect 5632 2261 5641 2295
rect 5641 2261 5675 2295
rect 5675 2261 5684 2295
rect 5632 2252 5684 2261
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 10508 2456 10560 2508
rect 12808 2431 12860 2440
rect 12808 2397 12817 2431
rect 12817 2397 12851 2431
rect 12851 2397 12860 2431
rect 12808 2388 12860 2397
rect 14372 2431 14424 2440
rect 14372 2397 14381 2431
rect 14381 2397 14415 2431
rect 14415 2397 14424 2431
rect 14372 2388 14424 2397
rect 13360 2320 13412 2372
rect 15476 2363 15528 2372
rect 15476 2329 15485 2363
rect 15485 2329 15519 2363
rect 15519 2329 15528 2363
rect 15476 2320 15528 2329
rect 15660 2363 15712 2372
rect 15660 2329 15669 2363
rect 15669 2329 15703 2363
rect 15703 2329 15712 2363
rect 15660 2320 15712 2329
rect 9588 2252 9640 2304
rect 6103 2150 6155 2202
rect 6167 2150 6219 2202
rect 6231 2150 6283 2202
rect 6295 2150 6347 2202
rect 11224 2150 11276 2202
rect 11288 2150 11340 2202
rect 11352 2150 11404 2202
rect 11416 2150 11468 2202
rect 1676 2048 1728 2100
rect 9496 2048 9548 2100
rect 4804 1980 4856 2032
rect 15660 1980 15712 2032
<< metal2 >>
rect 18 18928 74 19728
rect 2042 18928 2098 19728
rect 4066 18928 4122 19728
rect 5906 18928 5962 19728
rect 7930 18928 7986 19728
rect 9770 18928 9826 19728
rect 11794 18928 11850 19728
rect 13634 18928 13690 19728
rect 15658 18928 15714 19728
rect 17498 18928 17554 19728
rect 32 17338 60 18928
rect 20 17332 72 17338
rect 20 17274 72 17280
rect 1860 17264 1912 17270
rect 1858 17232 1860 17241
rect 1912 17232 1914 17241
rect 1676 17196 1728 17202
rect 1858 17167 1914 17176
rect 1676 17138 1728 17144
rect 1492 15700 1544 15706
rect 1492 15642 1544 15648
rect 1504 12782 1532 15642
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1596 13938 1624 14214
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1504 12238 1532 12718
rect 1688 12442 1716 17138
rect 2056 16522 2084 18928
rect 4080 17898 4108 18928
rect 4080 17870 4200 17898
rect 4172 17270 4200 17870
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 5920 17202 5948 18928
rect 6077 17436 6373 17456
rect 6133 17434 6157 17436
rect 6213 17434 6237 17436
rect 6293 17434 6317 17436
rect 6155 17382 6157 17434
rect 6219 17382 6231 17434
rect 6293 17382 6295 17434
rect 6133 17380 6157 17382
rect 6213 17380 6237 17382
rect 6293 17380 6317 17382
rect 6077 17360 6373 17380
rect 7944 17270 7972 18928
rect 9784 17338 9812 18928
rect 11198 17436 11494 17456
rect 11254 17434 11278 17436
rect 11334 17434 11358 17436
rect 11414 17434 11438 17436
rect 11276 17382 11278 17434
rect 11340 17382 11352 17434
rect 11414 17382 11416 17434
rect 11254 17380 11278 17382
rect 11334 17380 11358 17382
rect 11414 17380 11438 17382
rect 11198 17360 11494 17380
rect 11808 17354 11836 18928
rect 13648 17490 13676 18928
rect 13648 17462 13860 17490
rect 9772 17332 9824 17338
rect 11808 17326 11928 17354
rect 9772 17274 9824 17280
rect 11900 17270 11928 17326
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 3516 16892 3812 16912
rect 3572 16890 3596 16892
rect 3652 16890 3676 16892
rect 3732 16890 3756 16892
rect 3594 16838 3596 16890
rect 3658 16838 3670 16890
rect 3732 16838 3734 16890
rect 3572 16836 3596 16838
rect 3652 16836 3676 16838
rect 3732 16836 3756 16838
rect 3516 16816 3812 16836
rect 3056 16720 3108 16726
rect 3056 16662 3108 16668
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2044 16516 2096 16522
rect 2044 16458 2096 16464
rect 2516 16454 2544 16526
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2516 15910 2544 16390
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2516 15706 2544 15846
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2136 15632 2188 15638
rect 2136 15574 2188 15580
rect 2148 14890 2176 15574
rect 2792 15502 2820 16526
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2424 15026 2452 15302
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2136 14884 2188 14890
rect 2136 14826 2188 14832
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1964 14249 1992 14350
rect 1950 14240 2006 14249
rect 1950 14175 2006 14184
rect 2044 13728 2096 13734
rect 2044 13670 2096 13676
rect 2056 12850 2084 13670
rect 2148 13530 2176 14826
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2136 13524 2188 13530
rect 2136 13466 2188 13472
rect 2424 13326 2452 14010
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 2056 12730 2084 12786
rect 1964 12702 2084 12730
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1768 12368 1820 12374
rect 1768 12310 1820 12316
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1504 11150 1532 12174
rect 1780 11762 1808 12310
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 1872 11529 1900 12582
rect 1964 12442 1992 12702
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 2056 12238 2084 12582
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2044 12232 2096 12238
rect 1964 12192 2044 12220
rect 1858 11520 1914 11529
rect 1858 11455 1914 11464
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1596 6390 1624 6598
rect 1584 6384 1636 6390
rect 1584 6326 1636 6332
rect 1688 6322 1716 6598
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 5817 1440 6190
rect 1398 5808 1454 5817
rect 1398 5743 1454 5752
rect 1400 5568 1452 5574
rect 1400 5510 1452 5516
rect 1412 3126 1440 5510
rect 1780 5234 1808 11154
rect 1964 10742 1992 12192
rect 2044 12174 2096 12180
rect 2148 11830 2176 12242
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2136 11824 2188 11830
rect 2136 11766 2188 11772
rect 2148 11642 2176 11766
rect 2056 11614 2176 11642
rect 2056 11150 2084 11614
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2148 11218 2176 11494
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 2240 10674 2268 12174
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 1872 10062 1900 10406
rect 2240 10266 2268 10610
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2424 10130 2452 10610
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1964 9722 1992 10066
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1872 8498 1900 8842
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1872 7546 1900 8434
rect 1964 8430 1992 8842
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1596 4826 1624 4966
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1596 4078 1624 4762
rect 1688 4622 1716 4966
rect 1780 4622 1808 5170
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1688 4146 1716 4558
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1400 3120 1452 3126
rect 1596 3097 1624 3470
rect 1400 3062 1452 3068
rect 1582 3088 1638 3097
rect 1780 3058 1808 3878
rect 1872 3534 1900 5646
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1964 3602 1992 4558
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1582 3023 1638 3032
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1872 2854 1900 3470
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 2056 2514 2084 9862
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2148 9178 2176 9522
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2240 8634 2268 9522
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2424 7002 2452 8366
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2516 5817 2544 14758
rect 2792 14618 2820 15438
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2976 14414 3004 14758
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2976 13938 3004 14350
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2608 13530 2636 13670
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2884 11898 2912 13262
rect 3068 12918 3096 16662
rect 3700 16652 3752 16658
rect 3700 16594 3752 16600
rect 3712 16114 3740 16594
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 4080 16130 4108 16526
rect 3988 16114 4108 16130
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3976 16108 4108 16114
rect 4028 16102 4108 16108
rect 3976 16050 4028 16056
rect 4080 15978 4108 16102
rect 4068 15972 4120 15978
rect 4068 15914 4120 15920
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 3516 15804 3812 15824
rect 3572 15802 3596 15804
rect 3652 15802 3676 15804
rect 3732 15802 3756 15804
rect 3594 15750 3596 15802
rect 3658 15750 3670 15802
rect 3732 15750 3734 15802
rect 3572 15748 3596 15750
rect 3652 15748 3676 15750
rect 3732 15748 3756 15750
rect 3516 15728 3812 15748
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 3160 14414 3188 15370
rect 3344 15026 3372 15506
rect 3988 15162 4016 15846
rect 4160 15428 4212 15434
rect 4160 15370 4212 15376
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3516 14716 3812 14736
rect 3572 14714 3596 14716
rect 3652 14714 3676 14716
rect 3732 14714 3756 14716
rect 3594 14662 3596 14714
rect 3658 14662 3670 14714
rect 3732 14662 3734 14714
rect 3572 14660 3596 14662
rect 3652 14660 3676 14662
rect 3732 14660 3756 14662
rect 3516 14640 3812 14660
rect 4172 14618 4200 15370
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4172 14414 4200 14554
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 3160 12986 3188 14350
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3252 13326 3280 13806
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3056 12912 3108 12918
rect 3056 12854 3108 12860
rect 3436 12850 3464 13874
rect 3804 13716 3832 13874
rect 3804 13688 3924 13716
rect 3516 13628 3812 13648
rect 3572 13626 3596 13628
rect 3652 13626 3676 13628
rect 3732 13626 3756 13628
rect 3594 13574 3596 13626
rect 3658 13574 3670 13626
rect 3732 13574 3734 13626
rect 3572 13572 3596 13574
rect 3652 13572 3676 13574
rect 3732 13572 3756 13574
rect 3516 13552 3812 13572
rect 3896 13530 3924 13688
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3896 12850 3924 13466
rect 3988 13326 4016 13874
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 13326 4108 13670
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3516 12540 3812 12560
rect 3572 12538 3596 12540
rect 3652 12538 3676 12540
rect 3732 12538 3756 12540
rect 3594 12486 3596 12538
rect 3658 12486 3670 12538
rect 3732 12486 3734 12538
rect 3572 12484 3596 12486
rect 3652 12484 3676 12486
rect 3732 12484 3756 12486
rect 3516 12464 3812 12484
rect 3988 11898 4016 13262
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 4080 12442 4108 12854
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2792 11014 2820 11562
rect 2884 11150 2912 11562
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2792 10810 2820 10950
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2884 10198 2912 10950
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2976 9450 3004 11630
rect 3436 11354 3464 11630
rect 3516 11452 3812 11472
rect 3572 11450 3596 11452
rect 3652 11450 3676 11452
rect 3732 11450 3756 11452
rect 3594 11398 3596 11450
rect 3658 11398 3670 11450
rect 3732 11398 3734 11450
rect 3572 11396 3596 11398
rect 3652 11396 3676 11398
rect 3732 11396 3756 11398
rect 3516 11376 3812 11396
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3896 10810 3924 11154
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3252 10062 3280 10542
rect 3516 10364 3812 10384
rect 3572 10362 3596 10364
rect 3652 10362 3676 10364
rect 3732 10362 3756 10364
rect 3594 10310 3596 10362
rect 3658 10310 3670 10362
rect 3732 10310 3734 10362
rect 3572 10308 3596 10310
rect 3652 10308 3676 10310
rect 3732 10308 3756 10310
rect 3516 10288 3812 10308
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 8537 2912 8774
rect 3068 8634 3096 9998
rect 3252 9926 3280 9998
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3252 9586 3280 9862
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3516 9276 3812 9296
rect 3572 9274 3596 9276
rect 3652 9274 3676 9276
rect 3732 9274 3756 9276
rect 3594 9222 3596 9274
rect 3658 9222 3670 9274
rect 3732 9222 3734 9274
rect 3572 9220 3596 9222
rect 3652 9220 3676 9222
rect 3732 9220 3756 9222
rect 3516 9200 3812 9220
rect 4080 9178 4108 11086
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2870 8528 2926 8537
rect 2596 8492 2648 8498
rect 2870 8463 2926 8472
rect 2596 8434 2648 8440
rect 2608 8090 2636 8434
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2608 7410 2636 8026
rect 2700 7478 2728 8366
rect 3516 8188 3812 8208
rect 3572 8186 3596 8188
rect 3652 8186 3676 8188
rect 3732 8186 3756 8188
rect 3594 8134 3596 8186
rect 3658 8134 3670 8186
rect 3732 8134 3734 8186
rect 3572 8132 3596 8134
rect 3652 8132 3676 8134
rect 3732 8132 3756 8134
rect 3516 8112 3812 8132
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 2792 7410 2820 7686
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2792 7002 2820 7346
rect 2884 7342 2912 7822
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 3516 7100 3812 7120
rect 3572 7098 3596 7100
rect 3652 7098 3676 7100
rect 3732 7098 3756 7100
rect 3594 7046 3596 7098
rect 3658 7046 3670 7098
rect 3732 7046 3734 7098
rect 3572 7044 3596 7046
rect 3652 7044 3676 7046
rect 3732 7044 3756 7046
rect 3516 7024 3812 7044
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 2792 5817 2820 6122
rect 2502 5808 2558 5817
rect 2502 5743 2558 5752
rect 2778 5808 2834 5817
rect 2778 5743 2834 5752
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2148 2990 2176 5510
rect 2792 5370 2820 5646
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2332 4554 2360 5170
rect 2884 5114 2912 6666
rect 3068 5846 3096 6666
rect 3252 6458 3280 6734
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3252 5846 3280 6394
rect 3792 6248 3844 6254
rect 3844 6196 3924 6202
rect 3792 6190 3924 6196
rect 3804 6174 3924 6190
rect 3516 6012 3812 6032
rect 3572 6010 3596 6012
rect 3652 6010 3676 6012
rect 3732 6010 3756 6012
rect 3594 5958 3596 6010
rect 3658 5958 3670 6010
rect 3732 5958 3734 6010
rect 3572 5956 3596 5958
rect 3652 5956 3676 5958
rect 3732 5956 3756 5958
rect 3516 5936 3812 5956
rect 3896 5914 3924 6174
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3056 5840 3108 5846
rect 3056 5782 3108 5788
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 2792 5086 2912 5114
rect 2320 4548 2372 4554
rect 2320 4490 2372 4496
rect 2332 3602 2360 4490
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2686 3496 2742 3505
rect 2686 3431 2742 3440
rect 2594 3224 2650 3233
rect 2594 3159 2596 3168
rect 2648 3159 2650 3168
rect 2596 3130 2648 3136
rect 2700 3058 2728 3431
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2792 2825 2820 5086
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2884 4146 2912 4966
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2778 2816 2834 2825
rect 2778 2751 2834 2760
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 2976 2446 3004 4422
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3160 3058 3188 3538
rect 3344 3516 3372 5306
rect 3436 5234 3464 5510
rect 3988 5386 4016 7346
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 3896 5358 4016 5386
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3436 4690 3464 5170
rect 3516 4924 3812 4944
rect 3572 4922 3596 4924
rect 3652 4922 3676 4924
rect 3732 4922 3756 4924
rect 3594 4870 3596 4922
rect 3658 4870 3670 4922
rect 3732 4870 3734 4922
rect 3572 4868 3596 4870
rect 3652 4868 3676 4870
rect 3732 4868 3756 4870
rect 3516 4848 3812 4868
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3516 3836 3812 3856
rect 3572 3834 3596 3836
rect 3652 3834 3676 3836
rect 3732 3834 3756 3836
rect 3594 3782 3596 3834
rect 3658 3782 3670 3834
rect 3732 3782 3734 3834
rect 3572 3780 3596 3782
rect 3652 3780 3676 3782
rect 3732 3780 3756 3782
rect 3516 3760 3812 3780
rect 3896 3641 3924 5358
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 3988 4622 4016 5238
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 4080 4554 4108 5578
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 3882 3632 3938 3641
rect 3882 3567 3938 3576
rect 3884 3528 3936 3534
rect 3344 3488 3884 3516
rect 3344 3126 3372 3488
rect 3884 3470 3936 3476
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 3528 3058 3556 3334
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3896 2854 3924 3470
rect 4080 3398 4108 4490
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4080 3194 4108 3334
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4264 2922 4292 17138
rect 4896 17060 4948 17066
rect 4896 17002 4948 17008
rect 4908 16522 4936 17002
rect 5092 16794 5120 17138
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 5000 16114 5028 16526
rect 5368 16250 5396 16526
rect 5460 16454 5488 17138
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6104 16590 6132 16934
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5460 16250 5488 16390
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5644 16182 5672 16390
rect 5632 16176 5684 16182
rect 5632 16118 5684 16124
rect 5828 16114 5856 16526
rect 6077 16348 6373 16368
rect 6133 16346 6157 16348
rect 6213 16346 6237 16348
rect 6293 16346 6317 16348
rect 6155 16294 6157 16346
rect 6219 16294 6231 16346
rect 6293 16294 6295 16346
rect 6133 16292 6157 16294
rect 6213 16292 6237 16294
rect 6293 16292 6317 16294
rect 6077 16272 6373 16292
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6077 15260 6373 15280
rect 6133 15258 6157 15260
rect 6213 15258 6237 15260
rect 6293 15258 6317 15260
rect 6155 15206 6157 15258
rect 6219 15206 6231 15258
rect 6293 15206 6295 15258
rect 6133 15204 6157 15206
rect 6213 15204 6237 15206
rect 6293 15204 6317 15206
rect 6077 15184 6373 15204
rect 6472 15162 6500 16050
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 4448 14414 4476 14894
rect 4528 14884 4580 14890
rect 4528 14826 4580 14832
rect 4540 14414 4568 14826
rect 5000 14414 5028 14894
rect 5460 14618 5488 14894
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 5000 13530 5028 14350
rect 6077 14172 6373 14192
rect 6133 14170 6157 14172
rect 6213 14170 6237 14172
rect 6293 14170 6317 14172
rect 6155 14118 6157 14170
rect 6219 14118 6231 14170
rect 6293 14118 6295 14170
rect 6133 14116 6157 14118
rect 6213 14116 6237 14118
rect 6293 14116 6317 14118
rect 6077 14096 6373 14116
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 5092 13326 5120 13874
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5184 12866 5212 13670
rect 5276 13326 5304 13874
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5276 12986 5304 13262
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5184 12850 5304 12866
rect 5184 12844 5316 12850
rect 5184 12838 5264 12844
rect 5264 12786 5316 12792
rect 5368 12782 5396 13874
rect 5448 13252 5500 13258
rect 5448 13194 5500 13200
rect 5460 12986 5488 13194
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5184 11898 5212 12718
rect 5552 12170 5580 13942
rect 6077 13084 6373 13104
rect 6133 13082 6157 13084
rect 6213 13082 6237 13084
rect 6293 13082 6317 13084
rect 6155 13030 6157 13082
rect 6219 13030 6231 13082
rect 6293 13030 6295 13082
rect 6133 13028 6157 13030
rect 6213 13028 6237 13030
rect 6293 13028 6317 13030
rect 6077 13008 6373 13028
rect 6932 12434 6960 17070
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 7024 15978 7052 16526
rect 7116 16114 7144 16594
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 7380 15088 7432 15094
rect 7380 15030 7432 15036
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7300 14414 7328 14894
rect 7392 14414 7420 15030
rect 7484 14498 7512 17002
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7576 16046 7604 16390
rect 8128 16250 8156 16934
rect 8220 16794 8248 17138
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8312 16590 8340 17206
rect 13832 17202 13860 17462
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 8638 16892 8934 16912
rect 8694 16890 8718 16892
rect 8774 16890 8798 16892
rect 8854 16890 8878 16892
rect 8716 16838 8718 16890
rect 8780 16838 8792 16890
rect 8854 16838 8856 16890
rect 8694 16836 8718 16838
rect 8774 16836 8798 16838
rect 8854 16836 8878 16838
rect 8638 16816 8934 16836
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 8312 16182 8340 16390
rect 8300 16176 8352 16182
rect 8300 16118 8352 16124
rect 8404 16114 8432 16526
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7576 14618 7604 14962
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7484 14470 7604 14498
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 13870 7236 14214
rect 7300 14074 7328 14350
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7208 12918 7236 13126
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 6932 12406 7052 12434
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5632 11824 5684 11830
rect 5632 11766 5684 11772
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4540 10742 4568 11630
rect 4632 11082 4660 11630
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4632 10810 4660 11018
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4528 10736 4580 10742
rect 4528 10678 4580 10684
rect 4896 10668 4948 10674
rect 5448 10668 5500 10674
rect 4948 10628 5028 10656
rect 4896 10610 4948 10616
rect 5000 10588 5028 10628
rect 5448 10610 5500 10616
rect 5080 10600 5132 10606
rect 5000 10560 5080 10588
rect 5080 10542 5132 10548
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4356 7886 4384 8978
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4448 8362 4476 8842
rect 5092 8634 5120 10542
rect 5460 10266 5488 10610
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4448 7886 4476 8298
rect 4632 7954 4660 8434
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4632 7546 4660 7890
rect 4724 7886 4752 8366
rect 5354 7984 5410 7993
rect 5354 7919 5410 7928
rect 5368 7886 5396 7919
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4618 7440 4674 7449
rect 4618 7375 4620 7384
rect 4672 7375 4674 7384
rect 4620 7346 4672 7352
rect 4802 7304 4858 7313
rect 4802 7239 4804 7248
rect 4856 7239 4858 7248
rect 4804 7210 4856 7216
rect 5552 7154 5580 11222
rect 5644 10538 5672 11766
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5632 10532 5684 10538
rect 5632 10474 5684 10480
rect 5644 10062 5672 10474
rect 5736 10062 5764 11630
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5736 9382 5764 9998
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5828 9518 5856 9930
rect 5920 9654 5948 10066
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5816 9512 5868 9518
rect 6012 9466 6040 12106
rect 6077 11996 6373 12016
rect 6133 11994 6157 11996
rect 6213 11994 6237 11996
rect 6293 11994 6317 11996
rect 6155 11942 6157 11994
rect 6219 11942 6231 11994
rect 6293 11942 6295 11994
rect 6133 11940 6157 11942
rect 6213 11940 6237 11942
rect 6293 11940 6317 11942
rect 6077 11920 6373 11940
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6932 11218 6960 11698
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7024 11098 7052 12406
rect 7208 12238 7236 12854
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6932 11070 7052 11098
rect 7104 11076 7156 11082
rect 6077 10908 6373 10928
rect 6133 10906 6157 10908
rect 6213 10906 6237 10908
rect 6293 10906 6317 10908
rect 6155 10854 6157 10906
rect 6219 10854 6231 10906
rect 6293 10854 6295 10906
rect 6133 10852 6157 10854
rect 6213 10852 6237 10854
rect 6293 10852 6317 10854
rect 6077 10832 6373 10852
rect 6840 10198 6868 11018
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 6077 9820 6373 9840
rect 6133 9818 6157 9820
rect 6213 9818 6237 9820
rect 6293 9818 6317 9820
rect 6155 9766 6157 9818
rect 6219 9766 6231 9818
rect 6293 9766 6295 9818
rect 6133 9764 6157 9766
rect 6213 9764 6237 9766
rect 6293 9764 6317 9766
rect 6077 9744 6373 9764
rect 5816 9454 5868 9460
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5828 9110 5856 9454
rect 5920 9438 6040 9466
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5736 7342 5764 8366
rect 5828 7818 5856 8366
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5828 7274 5856 7754
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5552 7126 5856 7154
rect 5354 6896 5410 6905
rect 4528 6860 4580 6866
rect 5354 6831 5410 6840
rect 4528 6802 4580 6808
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4448 5914 4476 6190
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4540 5710 4568 6802
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 6458 4936 6734
rect 5368 6662 5396 6831
rect 5448 6792 5500 6798
rect 5500 6752 5672 6780
rect 5448 6734 5500 6740
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5460 6458 5488 6598
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 4908 6304 4936 6394
rect 4724 6276 4936 6304
rect 4724 5710 4752 6276
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5460 6118 5488 6190
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5460 5846 5488 6054
rect 5552 5914 5580 6190
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5092 5386 5120 5646
rect 4908 5358 5120 5386
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4356 4078 4384 4558
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4356 3670 4384 4014
rect 4540 3670 4568 4218
rect 4816 3942 4844 4694
rect 4908 4282 4936 5358
rect 5092 5302 5120 5358
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 5644 5234 5672 6752
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 5000 4622 5028 5034
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 5092 4622 5120 4966
rect 5184 4826 5212 5170
rect 5552 5114 5580 5170
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5460 5086 5580 5114
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5368 4622 5396 5034
rect 5460 4758 5488 5086
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4344 3664 4396 3670
rect 4344 3606 4396 3612
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4436 2984 4488 2990
rect 4434 2952 4436 2961
rect 4488 2952 4490 2961
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 4252 2916 4304 2922
rect 4434 2887 4490 2896
rect 4252 2858 4304 2864
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3516 2748 3812 2768
rect 3572 2746 3596 2748
rect 3652 2746 3676 2748
rect 3732 2746 3756 2748
rect 3594 2694 3596 2746
rect 3658 2694 3670 2746
rect 3732 2694 3734 2746
rect 3572 2692 3596 2694
rect 3652 2692 3676 2694
rect 3732 2692 3756 2694
rect 3516 2672 3812 2692
rect 4080 2446 4108 2858
rect 4724 2582 4752 3878
rect 5184 3534 5212 4422
rect 5368 4146 5396 4558
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 3194 5304 3402
rect 5460 3398 5488 4014
rect 5644 3618 5672 5170
rect 5736 4554 5764 5510
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5552 3590 5672 3618
rect 5724 3664 5776 3670
rect 5724 3606 5776 3612
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5552 3074 5580 3590
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5644 3233 5672 3470
rect 5630 3224 5686 3233
rect 5630 3159 5686 3168
rect 5460 3046 5580 3074
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 32 800 60 2382
rect 1688 2106 1716 2382
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 3884 2372 3936 2378
rect 3884 2314 3936 2320
rect 1676 2100 1728 2106
rect 1676 2042 1728 2048
rect 1872 800 1900 2314
rect 3896 800 3924 2314
rect 4816 2038 4844 2450
rect 5460 2446 5488 3046
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5552 2378 5580 2926
rect 5736 2666 5764 3606
rect 5644 2638 5764 2666
rect 5644 2514 5672 2638
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5828 2446 5856 7126
rect 5920 6798 5948 9438
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6012 8566 6040 9318
rect 6077 8732 6373 8752
rect 6133 8730 6157 8732
rect 6213 8730 6237 8732
rect 6293 8730 6317 8732
rect 6155 8678 6157 8730
rect 6219 8678 6231 8730
rect 6293 8678 6295 8730
rect 6133 8676 6157 8678
rect 6213 8676 6237 8678
rect 6293 8676 6317 8678
rect 6077 8656 6373 8676
rect 6932 8566 6960 11070
rect 7104 11018 7156 11024
rect 7116 10674 7144 11018
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7116 10266 7144 10610
rect 7208 10470 7236 11698
rect 7300 10690 7328 12378
rect 7484 12238 7512 12582
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7392 11218 7420 11630
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7380 11076 7432 11082
rect 7484 11064 7512 11698
rect 7576 11082 7604 14470
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 8036 14074 8064 14350
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7668 12306 7696 12786
rect 7852 12442 7880 13194
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7656 12300 7708 12306
rect 7944 12288 7972 13874
rect 7656 12242 7708 12248
rect 7760 12260 7972 12288
rect 7668 11898 7696 12242
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7432 11036 7512 11064
rect 7564 11076 7616 11082
rect 7380 11018 7432 11024
rect 7564 11018 7616 11024
rect 7392 10810 7420 11018
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7484 10690 7512 10746
rect 7300 10662 7512 10690
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7012 9716 7064 9722
rect 7392 9674 7420 10542
rect 7484 9994 7512 10662
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7012 9658 7064 9664
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6077 7644 6373 7664
rect 6133 7642 6157 7644
rect 6213 7642 6237 7644
rect 6293 7642 6317 7644
rect 6155 7590 6157 7642
rect 6219 7590 6231 7642
rect 6293 7590 6295 7642
rect 6133 7588 6157 7590
rect 6213 7588 6237 7590
rect 6293 7588 6317 7590
rect 6077 7568 6373 7588
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5920 5953 5948 6734
rect 6077 6556 6373 6576
rect 6133 6554 6157 6556
rect 6213 6554 6237 6556
rect 6293 6554 6317 6556
rect 6155 6502 6157 6554
rect 6219 6502 6231 6554
rect 6293 6502 6295 6554
rect 6133 6500 6157 6502
rect 6213 6500 6237 6502
rect 6293 6500 6317 6502
rect 6077 6480 6373 6500
rect 6472 6361 6500 8230
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6564 7857 6592 8026
rect 7024 7936 7052 9658
rect 7208 9646 7420 9674
rect 7208 9450 7236 9646
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 6840 7908 7052 7936
rect 6644 7880 6696 7886
rect 6550 7848 6606 7857
rect 6644 7822 6696 7828
rect 6550 7783 6606 7792
rect 6656 7721 6684 7822
rect 6736 7744 6788 7750
rect 6642 7712 6698 7721
rect 6736 7686 6788 7692
rect 6642 7647 6698 7656
rect 6748 7410 6776 7686
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6840 6882 6868 7908
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6748 6854 6868 6882
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6656 6633 6684 6734
rect 6642 6624 6698 6633
rect 6642 6559 6698 6568
rect 6458 6352 6514 6361
rect 6458 6287 6514 6296
rect 6552 6316 6604 6322
rect 5906 5944 5962 5953
rect 5906 5879 5962 5888
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5920 4622 5948 5646
rect 6472 5642 6500 6287
rect 6552 6258 6604 6264
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6564 5574 6592 6258
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6077 5468 6373 5488
rect 6133 5466 6157 5468
rect 6213 5466 6237 5468
rect 6293 5466 6317 5468
rect 6155 5414 6157 5466
rect 6219 5414 6231 5466
rect 6293 5414 6295 5466
rect 6133 5412 6157 5414
rect 6213 5412 6237 5414
rect 6293 5412 6317 5414
rect 6077 5392 6373 5412
rect 6656 5166 6684 6190
rect 6748 5794 6776 6854
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6840 6322 6868 6734
rect 6932 6610 6960 7482
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7024 7041 7052 7278
rect 7116 7274 7144 7686
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7010 7032 7066 7041
rect 7010 6967 7066 6976
rect 7116 6866 7144 7210
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7208 6780 7236 9386
rect 7300 7886 7328 9522
rect 7484 9466 7512 9930
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7576 9586 7604 9862
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7392 9438 7512 9466
rect 7392 8514 7420 9438
rect 7576 9042 7604 9522
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7484 8634 7512 8910
rect 7564 8900 7616 8906
rect 7668 8888 7696 10950
rect 7760 10606 7788 12260
rect 8220 12186 8248 15846
rect 8638 15804 8934 15824
rect 8694 15802 8718 15804
rect 8774 15802 8798 15804
rect 8854 15802 8878 15804
rect 8716 15750 8718 15802
rect 8780 15750 8792 15802
rect 8854 15750 8856 15802
rect 8694 15748 8718 15750
rect 8774 15748 8798 15750
rect 8854 15748 8878 15750
rect 8638 15728 8934 15748
rect 9232 15502 9260 16458
rect 9324 16250 9352 17070
rect 9416 16590 9444 17138
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10244 16590 10272 16934
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 10336 16114 10364 17138
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10428 16250 10456 16594
rect 11532 16522 11560 16934
rect 11520 16516 11572 16522
rect 11520 16458 11572 16464
rect 11198 16348 11494 16368
rect 11254 16346 11278 16348
rect 11334 16346 11358 16348
rect 11414 16346 11438 16348
rect 11276 16294 11278 16346
rect 11340 16294 11352 16346
rect 11414 16294 11416 16346
rect 11254 16292 11278 16294
rect 11334 16292 11358 16294
rect 11414 16292 11438 16294
rect 11198 16272 11494 16292
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10336 15706 10364 16050
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10888 15502 10916 15914
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 11072 15434 11100 16118
rect 11716 16046 11744 17138
rect 11808 16794 11836 17138
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11808 16114 11836 16730
rect 11900 16590 11928 16934
rect 12084 16658 12112 17138
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8496 14618 8524 14894
rect 8638 14716 8934 14736
rect 8694 14714 8718 14716
rect 8774 14714 8798 14716
rect 8854 14714 8878 14716
rect 8716 14662 8718 14714
rect 8780 14662 8792 14714
rect 8854 14662 8856 14714
rect 8694 14660 8718 14662
rect 8774 14660 8798 14662
rect 8854 14660 8878 14662
rect 8638 14640 8934 14660
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 8312 13870 8340 14350
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8312 13530 8340 13806
rect 8638 13628 8934 13648
rect 8694 13626 8718 13628
rect 8774 13626 8798 13628
rect 8854 13626 8878 13628
rect 8716 13574 8718 13626
rect 8780 13574 8792 13626
rect 8854 13574 8856 13626
rect 8694 13572 8718 13574
rect 8774 13572 8798 13574
rect 8854 13572 8878 13574
rect 8638 13552 8934 13572
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 9140 13326 9168 14350
rect 9232 13734 9260 14350
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9232 13326 9260 13670
rect 9508 13326 9536 13806
rect 9600 13462 9628 13874
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 8772 12850 8800 13262
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8956 12986 8984 13126
rect 9140 12986 9168 13262
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8312 12306 8340 12718
rect 9324 12646 9352 12854
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 8638 12540 8934 12560
rect 8694 12538 8718 12540
rect 8774 12538 8798 12540
rect 8854 12538 8878 12540
rect 8716 12486 8718 12538
rect 8780 12486 8792 12538
rect 8854 12486 8856 12538
rect 8694 12484 8718 12486
rect 8774 12484 8798 12486
rect 8854 12484 8878 12486
rect 8638 12464 8934 12484
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 7852 12158 8248 12186
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7760 9994 7788 10406
rect 7748 9988 7800 9994
rect 7748 9930 7800 9936
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7760 8906 7788 9522
rect 7616 8860 7696 8888
rect 7564 8842 7616 8848
rect 7668 8786 7696 8860
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 7668 8758 7788 8786
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7392 8486 7604 8514
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7392 8090 7420 8366
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7208 6752 7328 6780
rect 7300 6662 7328 6752
rect 7288 6656 7340 6662
rect 6932 6582 7236 6610
rect 7288 6598 7340 6604
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 7024 5846 7052 6190
rect 7012 5840 7064 5846
rect 6748 5766 6868 5794
rect 7012 5782 7064 5788
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6748 5370 6776 5646
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6840 5098 6868 5766
rect 7024 5234 7052 5782
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 6077 4380 6373 4400
rect 6133 4378 6157 4380
rect 6213 4378 6237 4380
rect 6293 4378 6317 4380
rect 6155 4326 6157 4378
rect 6219 4326 6231 4378
rect 6293 4326 6295 4378
rect 6133 4324 6157 4326
rect 6213 4324 6237 4326
rect 6293 4324 6317 4326
rect 6077 4304 6373 4324
rect 6932 4146 6960 5170
rect 7208 4622 7236 6582
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7208 4146 7236 4558
rect 7300 4321 7328 6598
rect 7286 4312 7342 4321
rect 7286 4247 7342 4256
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 5920 3534 5948 3606
rect 6104 3534 6132 3946
rect 6748 3534 6776 4082
rect 6828 4072 6880 4078
rect 7116 4049 7144 4082
rect 6828 4014 6880 4020
rect 7102 4040 7158 4049
rect 5908 3528 5960 3534
rect 6092 3528 6144 3534
rect 5908 3470 5960 3476
rect 6090 3496 6092 3505
rect 6736 3528 6788 3534
rect 6144 3496 6146 3505
rect 6736 3470 6788 3476
rect 6090 3431 6146 3440
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5920 2650 5948 2994
rect 6012 2990 6040 3334
rect 6077 3292 6373 3312
rect 6133 3290 6157 3292
rect 6213 3290 6237 3292
rect 6293 3290 6317 3292
rect 6155 3238 6157 3290
rect 6219 3238 6231 3290
rect 6293 3238 6295 3290
rect 6133 3236 6157 3238
rect 6213 3236 6237 3238
rect 6293 3236 6317 3238
rect 6077 3216 6373 3236
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6564 2514 6592 3334
rect 6748 3074 6776 3470
rect 6840 3466 6868 4014
rect 6920 4004 6972 4010
rect 7102 3975 7158 3984
rect 6920 3946 6972 3952
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6748 3046 6868 3074
rect 6840 2990 6868 3046
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6748 2446 6776 2926
rect 6932 2650 6960 3946
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7116 3097 7144 3674
rect 7194 3496 7250 3505
rect 7194 3431 7196 3440
rect 7248 3431 7250 3440
rect 7196 3402 7248 3408
rect 7288 3120 7340 3126
rect 7102 3088 7158 3097
rect 7102 3023 7158 3032
rect 7286 3088 7288 3097
rect 7340 3088 7342 3097
rect 7286 3023 7342 3032
rect 7116 2990 7144 3023
rect 7104 2984 7156 2990
rect 7010 2952 7066 2961
rect 7104 2926 7156 2932
rect 7010 2887 7012 2896
rect 7064 2887 7066 2896
rect 7012 2858 7064 2864
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 7116 2378 7144 2790
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 4804 2032 4856 2038
rect 4804 1974 4856 1980
rect 5644 1170 5672 2246
rect 6077 2204 6373 2224
rect 6133 2202 6157 2204
rect 6213 2202 6237 2204
rect 6293 2202 6317 2204
rect 6155 2150 6157 2202
rect 6219 2150 6231 2202
rect 6293 2150 6295 2202
rect 6133 2148 6157 2150
rect 6213 2148 6237 2150
rect 6293 2148 6317 2150
rect 6077 2128 6373 2148
rect 5644 1142 5764 1170
rect 5736 800 5764 1142
rect 18 0 74 800
rect 1858 0 1914 800
rect 3882 0 3938 800
rect 5722 0 5778 800
rect 7392 762 7420 7890
rect 7576 7818 7604 8486
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7470 7576 7526 7585
rect 7470 7511 7472 7520
rect 7524 7511 7526 7520
rect 7472 7482 7524 7488
rect 7760 7478 7788 8758
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7472 7404 7524 7410
rect 7656 7404 7708 7410
rect 7524 7364 7604 7392
rect 7472 7346 7524 7352
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7484 7002 7512 7142
rect 7576 7002 7604 7364
rect 7656 7346 7708 7352
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7472 6792 7524 6798
rect 7470 6760 7472 6769
rect 7524 6760 7526 6769
rect 7470 6695 7526 6704
rect 7668 6662 7696 7346
rect 7656 6656 7708 6662
rect 7654 6624 7656 6633
rect 7708 6624 7710 6633
rect 7654 6559 7710 6568
rect 7760 5930 7788 7414
rect 7852 6497 7880 12158
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7944 10062 7972 11766
rect 8036 11286 8064 12038
rect 8404 11830 8432 12038
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 8036 10130 8064 11222
rect 8128 10606 8156 11562
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 11354 8432 11494
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8496 11150 8524 11562
rect 8638 11452 8934 11472
rect 8694 11450 8718 11452
rect 8774 11450 8798 11452
rect 8854 11450 8878 11452
rect 8716 11398 8718 11450
rect 8780 11398 8792 11450
rect 8854 11398 8856 11450
rect 8694 11396 8718 11398
rect 8774 11396 8798 11398
rect 8854 11396 8878 11398
rect 8638 11376 8934 11396
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8220 10810 8248 10950
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8404 10674 8432 10950
rect 9416 10742 9444 13194
rect 9508 12646 9536 13262
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9692 12238 9720 12786
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9876 12238 9904 12718
rect 10152 12434 10180 14214
rect 10336 13326 10364 15302
rect 11198 15260 11494 15280
rect 11254 15258 11278 15260
rect 11334 15258 11358 15260
rect 11414 15258 11438 15260
rect 11276 15206 11278 15258
rect 11340 15206 11352 15258
rect 11414 15206 11416 15258
rect 11254 15204 11278 15206
rect 11334 15204 11358 15206
rect 11414 15204 11438 15206
rect 11198 15184 11494 15204
rect 11900 15162 11928 16526
rect 12176 16454 12204 17138
rect 12900 17060 12952 17066
rect 12900 17002 12952 17008
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12728 16574 12756 16934
rect 12728 16546 12848 16574
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 12268 15502 12296 15982
rect 12532 15632 12584 15638
rect 12532 15574 12584 15580
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 11348 14618 11376 14962
rect 11624 14958 11652 15030
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10980 14074 11008 14418
rect 11624 14414 11652 14894
rect 11992 14618 12020 14894
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11198 14172 11494 14192
rect 11254 14170 11278 14172
rect 11334 14170 11358 14172
rect 11414 14170 11438 14172
rect 11276 14118 11278 14170
rect 11340 14118 11352 14170
rect 11414 14118 11416 14170
rect 11254 14116 11278 14118
rect 11334 14116 11358 14118
rect 11414 14116 11438 14118
rect 11198 14096 11494 14116
rect 11624 14074 11652 14350
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 10980 13512 11008 14010
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11060 13524 11112 13530
rect 10888 13484 11060 13512
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10152 12406 10272 12434
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9692 11898 9720 12174
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9784 11830 9812 12106
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9508 11354 9536 11698
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9404 10736 9456 10742
rect 9404 10678 9456 10684
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 7944 6769 7972 7346
rect 8036 7177 8064 10066
rect 8128 9722 8156 10542
rect 8404 10062 8432 10610
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8638 10364 8934 10384
rect 8694 10362 8718 10364
rect 8774 10362 8798 10364
rect 8854 10362 8878 10364
rect 8716 10310 8718 10362
rect 8780 10310 8792 10362
rect 8854 10310 8856 10362
rect 8694 10308 8718 10310
rect 8774 10308 8798 10310
rect 8854 10308 8878 10310
rect 8638 10288 8934 10308
rect 9048 10062 9076 10406
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8312 8974 8340 9386
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 8786 8340 8910
rect 8220 8758 8340 8786
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8128 7886 8156 8434
rect 8220 8022 8248 8758
rect 8404 8430 8432 9454
rect 8638 9276 8934 9296
rect 8694 9274 8718 9276
rect 8774 9274 8798 9276
rect 8854 9274 8878 9276
rect 8716 9222 8718 9274
rect 8780 9222 8792 9274
rect 8854 9222 8856 9274
rect 8694 9220 8718 9222
rect 8774 9220 8798 9222
rect 8854 9220 8878 9222
rect 8638 9200 8934 9220
rect 9048 8922 9076 9998
rect 9140 9926 9168 10542
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9140 9042 9168 9862
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9048 8894 9168 8922
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7206 8156 7822
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8116 7200 8168 7206
rect 8022 7168 8078 7177
rect 8116 7142 8168 7148
rect 8022 7103 8078 7112
rect 8036 6934 8064 7103
rect 8024 6928 8076 6934
rect 8024 6870 8076 6876
rect 8220 6882 8248 7754
rect 8312 7698 8340 8298
rect 8404 8090 8432 8366
rect 8638 8188 8934 8208
rect 8694 8186 8718 8188
rect 8774 8186 8798 8188
rect 8854 8186 8878 8188
rect 8716 8134 8718 8186
rect 8780 8134 8792 8186
rect 8854 8134 8856 8186
rect 8694 8132 8718 8134
rect 8774 8132 8798 8134
rect 8854 8132 8878 8134
rect 8638 8112 8934 8132
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 9048 8022 9076 8434
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 8390 7712 8446 7721
rect 8312 7670 8390 7698
rect 8390 7647 8446 7656
rect 8298 7576 8354 7585
rect 8404 7546 8432 7647
rect 8298 7511 8354 7520
rect 8392 7540 8444 7546
rect 8312 7342 8340 7511
rect 8392 7482 8444 7488
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8404 6882 8432 7482
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8496 7177 8524 7346
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 8482 7168 8538 7177
rect 8482 7103 8538 7112
rect 8638 7100 8934 7120
rect 8694 7098 8718 7100
rect 8774 7098 8798 7100
rect 8854 7098 8878 7100
rect 8716 7046 8718 7098
rect 8780 7046 8792 7098
rect 8854 7046 8856 7098
rect 8694 7044 8718 7046
rect 8774 7044 8798 7046
rect 8854 7044 8878 7046
rect 8482 7032 8538 7041
rect 8638 7024 8934 7044
rect 9048 6984 9076 7210
rect 8538 6976 9076 6984
rect 8482 6967 9076 6976
rect 8496 6956 9076 6967
rect 9140 6905 9168 8894
rect 9416 7818 9444 10678
rect 9508 10674 9536 11086
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 10674 9720 11018
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9508 9722 9536 10610
rect 9692 10198 9720 10610
rect 9784 10266 9812 11766
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9876 9994 9904 11086
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 10060 10674 10088 10950
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 10266 9996 10542
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9600 8974 9628 9522
rect 9692 9382 9720 9862
rect 9876 9738 9904 9930
rect 9784 9722 9904 9738
rect 9968 9722 9996 10202
rect 10152 9926 10180 10406
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 9772 9716 9904 9722
rect 9824 9710 9904 9716
rect 9956 9716 10008 9722
rect 9772 9658 9824 9664
rect 9956 9658 10008 9664
rect 9956 9604 10008 9610
rect 9956 9546 10008 9552
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9126 6896 9182 6905
rect 8220 6854 8340 6882
rect 8404 6854 8524 6882
rect 8208 6792 8260 6798
rect 7930 6760 7986 6769
rect 8208 6734 8260 6740
rect 7930 6695 7986 6704
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 7838 6488 7894 6497
rect 7838 6423 7894 6432
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 7576 5902 7788 5930
rect 7576 5710 7604 5902
rect 7656 5840 7708 5846
rect 7656 5782 7708 5788
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7484 5234 7512 5578
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7484 2650 7512 5170
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7576 2446 7604 5306
rect 7668 5166 7696 5782
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7760 4078 7788 5902
rect 7852 5234 7880 6258
rect 7944 5778 7972 6394
rect 8036 6322 8064 6598
rect 8220 6458 8248 6734
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8312 6338 8340 6854
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8220 6310 8340 6338
rect 8404 6322 8432 6734
rect 8392 6316 8444 6322
rect 8220 6202 8248 6310
rect 8392 6258 8444 6264
rect 8496 6254 8524 6854
rect 8760 6860 8812 6866
rect 9416 6866 9444 7754
rect 9126 6831 9182 6840
rect 9404 6860 9456 6866
rect 8760 6802 8812 6808
rect 9404 6802 9456 6808
rect 8772 6458 8800 6802
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8036 6174 8248 6202
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7852 4826 7880 5170
rect 8036 5030 8064 6174
rect 8312 6100 8340 6190
rect 8128 6072 8340 6100
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 8036 4282 8064 4966
rect 8128 4486 8156 6072
rect 8638 6012 8934 6032
rect 8694 6010 8718 6012
rect 8774 6010 8798 6012
rect 8854 6010 8878 6012
rect 8716 5958 8718 6010
rect 8780 5958 8792 6010
rect 8854 5958 8856 6010
rect 8694 5956 8718 5958
rect 8774 5956 8798 5958
rect 8854 5956 8878 5958
rect 8206 5944 8262 5953
rect 8638 5936 8934 5956
rect 8206 5879 8262 5888
rect 8220 5846 8248 5879
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8220 5370 8248 5510
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8312 5166 8340 5646
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7840 4208 7892 4214
rect 8220 4185 8248 5034
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4622 8340 4966
rect 8404 4826 8432 5646
rect 8484 5636 8536 5642
rect 8484 5578 8536 5584
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8390 4312 8446 4321
rect 8390 4247 8446 4256
rect 7840 4150 7892 4156
rect 8206 4176 8262 4185
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7746 3632 7802 3641
rect 7746 3567 7802 3576
rect 7760 2922 7788 3567
rect 7852 3058 7880 4150
rect 8206 4111 8262 4120
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 8036 3670 8064 3878
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 8036 2446 8064 3606
rect 8220 3534 8248 4111
rect 8298 4040 8354 4049
rect 8298 3975 8354 3984
rect 8312 3738 8340 3975
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8298 3496 8354 3505
rect 8298 3431 8354 3440
rect 8312 2650 8340 3431
rect 8404 3398 8432 4247
rect 8496 4010 8524 5578
rect 8638 4924 8934 4944
rect 8694 4922 8718 4924
rect 8774 4922 8798 4924
rect 8854 4922 8878 4924
rect 8716 4870 8718 4922
rect 8780 4870 8792 4922
rect 8854 4870 8856 4922
rect 8694 4868 8718 4870
rect 8774 4868 8798 4870
rect 8854 4868 8878 4870
rect 8638 4848 8934 4868
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 8956 4486 8984 4558
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 9232 4321 9260 4558
rect 9312 4548 9364 4554
rect 9312 4490 9364 4496
rect 9218 4312 9274 4321
rect 9218 4247 9274 4256
rect 9220 4208 9272 4214
rect 9220 4150 9272 4156
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8638 3836 8934 3856
rect 8694 3834 8718 3836
rect 8774 3834 8798 3836
rect 8854 3834 8878 3836
rect 8716 3782 8718 3834
rect 8780 3782 8792 3834
rect 8854 3782 8856 3834
rect 8694 3780 8718 3782
rect 8774 3780 8798 3782
rect 8854 3780 8878 3782
rect 8638 3760 8934 3780
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8496 3058 8524 3606
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8680 3058 8708 3470
rect 9140 3194 9168 3674
rect 9232 3534 9260 4150
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 8760 3120 8812 3126
rect 8758 3088 8760 3097
rect 8812 3088 8814 3097
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8668 3052 8720 3058
rect 8758 3023 8814 3032
rect 8668 2994 8720 3000
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8404 2530 8432 2858
rect 8638 2748 8934 2768
rect 8694 2746 8718 2748
rect 8774 2746 8798 2748
rect 8854 2746 8878 2748
rect 8716 2694 8718 2746
rect 8780 2694 8792 2746
rect 8854 2694 8856 2746
rect 8694 2692 8718 2694
rect 8774 2692 8798 2694
rect 8854 2692 8878 2694
rect 8638 2672 8934 2692
rect 8312 2514 8432 2530
rect 8300 2508 8432 2514
rect 8352 2502 8432 2508
rect 8300 2450 8352 2456
rect 9140 2446 9168 3130
rect 9232 2922 9260 3470
rect 9324 3398 9352 4490
rect 9402 4176 9458 4185
rect 9402 4111 9404 4120
rect 9456 4111 9458 4120
rect 9404 4082 9456 4088
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9508 3738 9536 4014
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 9416 2582 9444 3538
rect 9600 2774 9628 8910
rect 9968 8498 9996 9546
rect 10152 9042 10180 9862
rect 10244 9178 10272 12406
rect 10336 11762 10364 13262
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10704 12918 10732 13126
rect 10888 12986 10916 13484
rect 11060 13466 11112 13472
rect 11164 13394 11192 13806
rect 11624 13802 11652 13874
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11348 13326 11376 13670
rect 11808 13394 11836 13874
rect 11900 13734 11928 13942
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11060 13252 11112 13258
rect 10980 13212 11060 13240
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10612 11150 10640 12310
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 11218 10732 11630
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 10538 10364 10950
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10336 10130 10364 10474
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 10152 8090 10180 8978
rect 10336 8634 10364 10066
rect 10428 9674 10456 10746
rect 10428 9646 10548 9674
rect 10520 9382 10548 9646
rect 10612 9586 10640 11086
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10324 8628 10376 8634
rect 10376 8588 10456 8616
rect 10324 8570 10376 8576
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 9692 7886 9720 8026
rect 9680 7880 9732 7886
rect 10048 7880 10100 7886
rect 9680 7822 9732 7828
rect 9862 7848 9918 7857
rect 9692 7546 9720 7822
rect 10048 7822 10100 7828
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 9862 7783 9918 7792
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9678 6760 9734 6769
rect 9678 6695 9734 6704
rect 9692 6390 9720 6695
rect 9770 6488 9826 6497
rect 9770 6423 9826 6432
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9784 6322 9812 6423
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9770 6216 9826 6225
rect 9770 6151 9772 6160
rect 9824 6151 9826 6160
rect 9772 6122 9824 6128
rect 9876 5710 9904 7783
rect 10060 7410 10088 7822
rect 10152 7546 10180 7822
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10336 6497 10364 6802
rect 10138 6488 10194 6497
rect 10138 6423 10194 6432
rect 10322 6488 10378 6497
rect 10322 6423 10378 6432
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9876 5302 9904 5646
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 10152 4826 10180 6423
rect 10322 6352 10378 6361
rect 10322 6287 10378 6296
rect 10336 6254 10364 6287
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10428 5574 10456 8588
rect 10520 8498 10548 9318
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10520 7324 10548 8434
rect 10704 7954 10732 11154
rect 10980 10810 11008 13212
rect 11060 13194 11112 13200
rect 11198 13084 11494 13104
rect 11254 13082 11278 13084
rect 11334 13082 11358 13084
rect 11414 13082 11438 13084
rect 11276 13030 11278 13082
rect 11340 13030 11352 13082
rect 11414 13030 11416 13082
rect 11254 13028 11278 13030
rect 11334 13028 11358 13030
rect 11414 13028 11438 13030
rect 11198 13008 11494 13028
rect 11992 12986 12020 13874
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 12084 13530 12112 13670
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 11072 12238 11100 12854
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 11440 12442 11468 12786
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 11072 10674 11100 12174
rect 11440 12170 11468 12378
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11198 11996 11494 12016
rect 11254 11994 11278 11996
rect 11334 11994 11358 11996
rect 11414 11994 11438 11996
rect 11276 11942 11278 11994
rect 11340 11942 11352 11994
rect 11414 11942 11416 11994
rect 11254 11940 11278 11942
rect 11334 11940 11358 11942
rect 11414 11940 11438 11942
rect 11198 11920 11494 11940
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11198 10908 11494 10928
rect 11254 10906 11278 10908
rect 11334 10906 11358 10908
rect 11414 10906 11438 10908
rect 11276 10854 11278 10906
rect 11340 10854 11352 10906
rect 11414 10854 11416 10906
rect 11254 10852 11278 10854
rect 11334 10852 11358 10854
rect 11414 10852 11438 10854
rect 11198 10832 11494 10852
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10888 10266 10916 10542
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10796 10130 10824 10202
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11072 9178 11100 9930
rect 11198 9820 11494 9840
rect 11254 9818 11278 9820
rect 11334 9818 11358 9820
rect 11414 9818 11438 9820
rect 11276 9766 11278 9818
rect 11340 9766 11352 9818
rect 11414 9766 11416 9818
rect 11254 9764 11278 9766
rect 11334 9764 11358 9766
rect 11414 9764 11438 9766
rect 11198 9744 11494 9764
rect 11624 9738 11652 11698
rect 11808 11694 11836 12174
rect 11992 11762 12020 12242
rect 12084 12238 12112 12786
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12084 11778 12112 12174
rect 12176 11898 12204 13194
rect 12268 12442 12296 15438
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 12360 15162 12388 15370
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12452 14006 12480 14282
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12360 13530 12388 13738
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12452 13258 12480 13670
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12452 12238 12480 12786
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11980 11756 12032 11762
rect 12084 11750 12296 11778
rect 11980 11698 12032 11704
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11900 11286 11928 11698
rect 11992 11354 12020 11698
rect 12072 11620 12124 11626
rect 12072 11562 12124 11568
rect 12084 11354 12112 11562
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11888 11280 11940 11286
rect 11888 11222 11940 11228
rect 11900 10810 11928 11222
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11808 10470 11836 10678
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11624 9710 11744 9738
rect 11716 9654 11744 9710
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11624 9178 11652 9522
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11198 8732 11494 8752
rect 11254 8730 11278 8732
rect 11334 8730 11358 8732
rect 11414 8730 11438 8732
rect 11276 8678 11278 8730
rect 11340 8678 11352 8730
rect 11414 8678 11416 8730
rect 11254 8676 11278 8678
rect 11334 8676 11358 8678
rect 11414 8676 11438 8678
rect 11198 8656 11494 8676
rect 11532 8566 11560 8842
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10612 7478 10640 7686
rect 10600 7472 10652 7478
rect 10600 7414 10652 7420
rect 10520 7296 10640 7324
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10508 5568 10560 5574
rect 10612 5556 10640 7296
rect 10704 6934 10732 7890
rect 10888 7886 10916 8230
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10888 7410 10916 7822
rect 11612 7812 11664 7818
rect 11612 7754 11664 7760
rect 11198 7644 11494 7664
rect 11254 7642 11278 7644
rect 11334 7642 11358 7644
rect 11414 7642 11438 7644
rect 11276 7590 11278 7642
rect 11340 7590 11352 7642
rect 11414 7590 11416 7642
rect 11254 7588 11278 7590
rect 11334 7588 11358 7590
rect 11414 7588 11438 7590
rect 11198 7568 11494 7588
rect 11150 7440 11206 7449
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10968 7404 11020 7410
rect 11150 7375 11206 7384
rect 10968 7346 11020 7352
rect 10980 7290 11008 7346
rect 10888 7262 11008 7290
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10704 6390 10732 6870
rect 10888 6730 10916 7262
rect 10966 7032 11022 7041
rect 11072 7002 11100 7278
rect 10966 6967 11022 6976
rect 11060 6996 11112 7002
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10980 6662 11008 6967
rect 11060 6938 11112 6944
rect 11164 6746 11192 7375
rect 11518 7304 11574 7313
rect 11518 7239 11574 7248
rect 11426 6896 11482 6905
rect 11426 6831 11482 6840
rect 11072 6718 11192 6746
rect 11440 6730 11468 6831
rect 11428 6724 11480 6730
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10796 5914 10824 6258
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10560 5528 10640 5556
rect 10692 5568 10744 5574
rect 10508 5510 10560 5516
rect 10692 5510 10744 5516
rect 10428 5370 10456 5510
rect 10520 5370 10548 5510
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10612 4128 10640 5170
rect 10704 5166 10732 5510
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10796 4554 10824 5850
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10980 5098 11008 5578
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 11072 4978 11100 6718
rect 11428 6666 11480 6672
rect 11198 6556 11494 6576
rect 11254 6554 11278 6556
rect 11334 6554 11358 6556
rect 11414 6554 11438 6556
rect 11276 6502 11278 6554
rect 11340 6502 11352 6554
rect 11414 6502 11416 6554
rect 11254 6500 11278 6502
rect 11334 6500 11358 6502
rect 11414 6500 11438 6502
rect 11198 6480 11494 6500
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11532 6338 11560 7239
rect 11624 7206 11652 7754
rect 11716 7206 11744 9590
rect 11900 7818 11928 10610
rect 11992 10266 12020 11290
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 11992 9042 12020 9930
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11440 5692 11468 6326
rect 11532 6310 11652 6338
rect 11520 5704 11572 5710
rect 11440 5664 11520 5692
rect 11520 5646 11572 5652
rect 11198 5468 11494 5488
rect 11254 5466 11278 5468
rect 11334 5466 11358 5468
rect 11414 5466 11438 5468
rect 11276 5414 11278 5466
rect 11340 5414 11352 5466
rect 11414 5414 11416 5466
rect 11254 5412 11278 5414
rect 11334 5412 11358 5414
rect 11414 5412 11438 5414
rect 11198 5392 11494 5412
rect 11624 5166 11652 6310
rect 11716 5166 11744 7142
rect 11796 6792 11848 6798
rect 11794 6760 11796 6769
rect 11848 6760 11850 6769
rect 11794 6695 11850 6704
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 6361 11836 6598
rect 11794 6352 11850 6361
rect 11794 6287 11850 6296
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11612 5160 11664 5166
rect 11612 5102 11664 5108
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 10888 4622 10916 4966
rect 11072 4950 11652 4978
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 10784 4140 10836 4146
rect 10612 4100 10784 4128
rect 10784 4082 10836 4088
rect 10796 4010 10824 4082
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 11072 3942 11100 4490
rect 11198 4380 11494 4400
rect 11254 4378 11278 4380
rect 11334 4378 11358 4380
rect 11414 4378 11438 4380
rect 11276 4326 11278 4378
rect 11340 4326 11352 4378
rect 11414 4326 11416 4378
rect 11254 4324 11278 4326
rect 11334 4324 11358 4326
rect 11414 4324 11438 4326
rect 11198 4304 11494 4324
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 9692 3058 9720 3878
rect 10336 3670 10364 3878
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 11072 3058 11100 3878
rect 11164 3534 11192 3878
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11198 3292 11494 3312
rect 11254 3290 11278 3292
rect 11334 3290 11358 3292
rect 11414 3290 11438 3292
rect 11276 3238 11278 3290
rect 11340 3238 11352 3290
rect 11414 3238 11416 3290
rect 11254 3236 11278 3238
rect 11334 3236 11358 3238
rect 11414 3236 11438 3238
rect 11198 3216 11494 3236
rect 11532 3194 11560 3538
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 10046 2952 10102 2961
rect 9508 2746 9628 2774
rect 9404 2576 9456 2582
rect 9404 2518 9456 2524
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9416 2378 9444 2518
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 9508 2106 9536 2746
rect 9876 2650 9904 2926
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9968 2446 9996 2926
rect 10046 2887 10102 2896
rect 10060 2582 10088 2887
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 10520 2514 10548 2994
rect 10508 2508 10560 2514
rect 10508 2450 10560 2456
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9496 2100 9548 2106
rect 9496 2042 9548 2048
rect 7668 870 7788 898
rect 7668 762 7696 870
rect 7760 800 7788 870
rect 9600 800 9628 2246
rect 11198 2204 11494 2224
rect 11254 2202 11278 2204
rect 11334 2202 11358 2204
rect 11414 2202 11438 2204
rect 11276 2150 11278 2202
rect 11340 2150 11352 2202
rect 11414 2150 11416 2202
rect 11254 2148 11278 2150
rect 11334 2148 11358 2150
rect 11414 2148 11438 2150
rect 11198 2128 11494 2148
rect 11624 800 11652 4950
rect 11716 4826 11744 5102
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11808 4622 11836 5170
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11900 4434 11928 7754
rect 11992 7410 12020 8978
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12084 7410 12112 8366
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11992 5234 12020 7346
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12084 6458 12112 6938
rect 12176 6458 12204 7482
rect 12268 7410 12296 11750
rect 12452 11082 12480 12174
rect 12544 11257 12572 15574
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12636 12714 12664 14758
rect 12728 13734 12756 14962
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12728 12442 12756 13670
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12820 12288 12848 16546
rect 12912 14074 12940 17002
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 13759 16892 14055 16912
rect 13815 16890 13839 16892
rect 13895 16890 13919 16892
rect 13975 16890 13999 16892
rect 13837 16838 13839 16890
rect 13901 16838 13913 16890
rect 13975 16838 13977 16890
rect 13815 16836 13839 16838
rect 13895 16836 13919 16838
rect 13975 16836 13999 16838
rect 13759 16816 14055 16836
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13464 16522 13492 16662
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13452 16516 13504 16522
rect 13452 16458 13504 16464
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13188 15706 13216 15982
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 12912 13938 12940 14010
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 13004 12986 13032 15642
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12912 12434 12940 12786
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 12912 12406 13032 12434
rect 12820 12260 12940 12288
rect 12530 11248 12586 11257
rect 12530 11183 12586 11192
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12452 9994 12480 10610
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 12544 9738 12572 10950
rect 12636 10418 12664 11018
rect 12820 10606 12848 11086
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12636 10390 12848 10418
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12452 9710 12572 9738
rect 12452 9042 12480 9710
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12360 8090 12388 8842
rect 12452 8566 12480 8978
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12452 7750 12480 8502
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12176 5574 12204 6394
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 11980 5228 12032 5234
rect 12268 5216 12296 7346
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12360 5574 12388 6258
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12452 5370 12480 5578
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 11980 5170 12032 5176
rect 12176 5188 12296 5216
rect 12440 5228 12492 5234
rect 11992 4554 12020 5170
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 11900 4406 12020 4434
rect 11992 4146 12020 4406
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 11808 2650 11836 3606
rect 12176 3602 12204 5188
rect 12440 5170 12492 5176
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 12268 3058 12296 5034
rect 12452 4486 12480 5170
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12452 4282 12480 4422
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12544 4146 12572 9522
rect 12636 8498 12664 9930
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12728 8294 12756 9318
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12348 3528 12400 3534
rect 12452 3516 12480 4082
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12400 3488 12480 3516
rect 12348 3470 12400 3476
rect 12544 3126 12572 3878
rect 12636 3670 12664 7278
rect 12728 7041 12756 7346
rect 12714 7032 12770 7041
rect 12714 6967 12770 6976
rect 12820 6746 12848 10390
rect 12912 9586 12940 12260
rect 13004 11354 13032 12406
rect 13188 12238 13216 12650
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13004 9926 13032 10610
rect 13096 10198 13124 11698
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13096 10062 13124 10134
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12912 7818 12940 8434
rect 13004 8362 13032 9862
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 13096 8634 13124 9386
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 12992 8356 13044 8362
rect 12992 8298 13044 8304
rect 12990 7984 13046 7993
rect 12990 7919 13046 7928
rect 12900 7812 12952 7818
rect 12900 7754 12952 7760
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 6905 12940 7142
rect 12898 6896 12954 6905
rect 12898 6831 12954 6840
rect 12728 6718 12848 6746
rect 12728 4554 12756 6718
rect 13004 6474 13032 7919
rect 13096 7886 13124 8570
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13084 7744 13136 7750
rect 13188 7732 13216 8570
rect 13280 8430 13308 14350
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13372 12850 13400 13194
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13372 12306 13400 12786
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13372 11082 13400 11562
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13464 9450 13492 16458
rect 13556 14074 13584 16594
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 14384 16454 14412 16526
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14384 16182 14412 16390
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 14476 16114 14504 16526
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 13759 15804 14055 15824
rect 13815 15802 13839 15804
rect 13895 15802 13919 15804
rect 13975 15802 13999 15804
rect 13837 15750 13839 15802
rect 13901 15750 13913 15802
rect 13975 15750 13977 15802
rect 13815 15748 13839 15750
rect 13895 15748 13919 15750
rect 13975 15748 13999 15750
rect 13759 15728 14055 15748
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 14004 14952 14056 14958
rect 14108 14906 14136 15370
rect 14056 14900 14136 14906
rect 14004 14894 14136 14900
rect 14016 14878 14136 14894
rect 13759 14716 14055 14736
rect 13815 14714 13839 14716
rect 13895 14714 13919 14716
rect 13975 14714 13999 14716
rect 13837 14662 13839 14714
rect 13901 14662 13913 14714
rect 13975 14662 13977 14714
rect 13815 14660 13839 14662
rect 13895 14660 13919 14662
rect 13975 14660 13999 14662
rect 13759 14640 14055 14660
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13556 11898 13584 13194
rect 13648 12434 13676 13942
rect 13759 13628 14055 13648
rect 13815 13626 13839 13628
rect 13895 13626 13919 13628
rect 13975 13626 13999 13628
rect 13837 13574 13839 13626
rect 13901 13574 13913 13626
rect 13975 13574 13977 13626
rect 13815 13572 13839 13574
rect 13895 13572 13919 13574
rect 13975 13572 13999 13574
rect 13759 13552 14055 13572
rect 14108 13530 14136 14878
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14200 13938 14228 14418
rect 14568 14362 14596 16934
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15212 16114 15240 16458
rect 15304 16182 15332 16458
rect 15396 16250 15424 17138
rect 15672 16574 15700 18928
rect 17512 17270 17540 18928
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 15752 17060 15804 17066
rect 15752 17002 15804 17008
rect 15764 16969 15792 17002
rect 15750 16960 15806 16969
rect 15750 16895 15806 16904
rect 15488 16546 15700 16574
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 14476 14334 14596 14362
rect 14384 13938 14412 14282
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14200 13530 14228 13874
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14292 13258 14320 13806
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 13759 12540 14055 12560
rect 13815 12538 13839 12540
rect 13895 12538 13919 12540
rect 13975 12538 13999 12540
rect 13837 12486 13839 12538
rect 13901 12486 13913 12538
rect 13975 12486 13977 12538
rect 13815 12484 13839 12486
rect 13895 12484 13919 12486
rect 13975 12484 13999 12486
rect 13759 12464 14055 12484
rect 14200 12442 14228 12786
rect 14188 12436 14240 12442
rect 13648 12406 13768 12434
rect 13740 12238 13768 12406
rect 14188 12378 14240 12384
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13740 11762 13768 12174
rect 14200 11830 14228 12242
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 14004 11756 14056 11762
rect 14056 11716 14136 11744
rect 14004 11698 14056 11704
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 11354 13676 11494
rect 13759 11452 14055 11472
rect 13815 11450 13839 11452
rect 13895 11450 13919 11452
rect 13975 11450 13999 11452
rect 13837 11398 13839 11450
rect 13901 11398 13913 11450
rect 13975 11398 13977 11450
rect 13815 11396 13839 11398
rect 13895 11396 13919 11398
rect 13975 11396 13999 11398
rect 13759 11376 14055 11396
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13556 10538 13584 11290
rect 14108 11150 14136 11716
rect 14200 11218 14228 11766
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13759 10364 14055 10384
rect 13815 10362 13839 10364
rect 13895 10362 13919 10364
rect 13975 10362 13999 10364
rect 13837 10310 13839 10362
rect 13901 10310 13913 10362
rect 13975 10310 13977 10362
rect 13815 10308 13839 10310
rect 13895 10308 13919 10310
rect 13975 10308 13999 10310
rect 13759 10288 14055 10308
rect 14108 10062 14136 11086
rect 14292 10810 14320 13194
rect 14384 12986 14412 13874
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14384 12238 14412 12786
rect 14476 12374 14504 14334
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14464 12368 14516 12374
rect 14464 12310 14516 12316
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14384 10674 14412 12174
rect 14476 11694 14504 12174
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 13556 9178 13584 9522
rect 13759 9276 14055 9296
rect 13815 9274 13839 9276
rect 13895 9274 13919 9276
rect 13975 9274 13999 9276
rect 13837 9222 13839 9274
rect 13901 9222 13913 9274
rect 13975 9222 13977 9274
rect 13815 9220 13839 9222
rect 13895 9220 13919 9222
rect 13975 9220 13999 9222
rect 13759 9200 14055 9220
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13452 9104 13504 9110
rect 13504 9052 13584 9058
rect 13452 9046 13584 9052
rect 13464 9030 13584 9046
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 13464 8634 13492 8842
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13372 7954 13400 8298
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13136 7704 13216 7732
rect 13084 7686 13136 7692
rect 13096 6662 13124 7686
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 13188 6934 13216 7414
rect 13176 6928 13228 6934
rect 13176 6870 13228 6876
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13004 6446 13124 6474
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12820 5914 12848 6258
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12912 5370 12940 6326
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12912 4554 12940 5102
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12900 4548 12952 4554
rect 12900 4490 12952 4496
rect 12728 4214 12756 4490
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 13004 4146 13032 5510
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12728 3466 12756 4014
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 12728 2650 12756 3402
rect 12820 3398 12848 3674
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12808 3120 12860 3126
rect 12808 3062 12860 3068
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12820 2446 12848 3062
rect 12912 2990 12940 3946
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 13096 2774 13124 6446
rect 13188 6322 13216 6666
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13188 4826 13216 6258
rect 13280 5522 13308 7822
rect 13372 7206 13400 7890
rect 13464 7750 13492 8230
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 5846 13400 7142
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13464 5710 13492 7686
rect 13556 7018 13584 9030
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13648 8022 13676 8502
rect 13759 8188 14055 8208
rect 13815 8186 13839 8188
rect 13895 8186 13919 8188
rect 13975 8186 13999 8188
rect 13837 8134 13839 8186
rect 13901 8134 13913 8186
rect 13975 8134 13977 8186
rect 13815 8132 13839 8134
rect 13895 8132 13919 8134
rect 13975 8132 13999 8134
rect 13759 8112 14055 8132
rect 14108 8090 14136 8910
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 13832 7410 13860 7482
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13759 7100 14055 7120
rect 13815 7098 13839 7100
rect 13895 7098 13919 7100
rect 13975 7098 13999 7100
rect 13837 7046 13839 7098
rect 13901 7046 13913 7098
rect 13975 7046 13977 7098
rect 13815 7044 13839 7046
rect 13895 7044 13919 7046
rect 13975 7044 13999 7046
rect 13759 7024 14055 7044
rect 13556 6990 13676 7018
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13556 6322 13584 6802
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13280 5494 13492 5522
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13372 4826 13400 5102
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13280 3652 13308 4694
rect 13372 3754 13400 4762
rect 13464 4010 13492 5494
rect 13556 5370 13584 5578
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13556 4758 13584 5306
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13372 3726 13492 3754
rect 13556 3738 13584 4558
rect 13280 3624 13400 3652
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13188 2854 13216 3130
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13280 2854 13308 2994
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13004 2746 13124 2774
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 7392 734 7696 762
rect 7746 0 7802 800
rect 9586 0 9642 800
rect 11610 0 11666 800
rect 13004 762 13032 2746
rect 13372 2378 13400 3624
rect 13464 3126 13492 3726
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13648 3210 13676 6990
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13740 6225 13768 6258
rect 13726 6216 13782 6225
rect 13726 6151 13782 6160
rect 13759 6012 14055 6032
rect 13815 6010 13839 6012
rect 13895 6010 13919 6012
rect 13975 6010 13999 6012
rect 13837 5958 13839 6010
rect 13901 5958 13913 6010
rect 13975 5958 13977 6010
rect 13815 5956 13839 5958
rect 13895 5956 13919 5958
rect 13975 5956 13999 5958
rect 13759 5936 14055 5956
rect 14108 5794 14136 7482
rect 13924 5766 14136 5794
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13740 5250 13768 5646
rect 13924 5302 13952 5766
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 13912 5296 13964 5302
rect 13740 5234 13860 5250
rect 13912 5238 13964 5244
rect 13740 5228 13872 5234
rect 13740 5222 13820 5228
rect 13820 5170 13872 5176
rect 13759 4924 14055 4944
rect 13815 4922 13839 4924
rect 13895 4922 13919 4924
rect 13975 4922 13999 4924
rect 13837 4870 13839 4922
rect 13901 4870 13913 4922
rect 13975 4870 13977 4922
rect 13815 4868 13839 4870
rect 13895 4868 13919 4870
rect 13975 4868 13999 4870
rect 13759 4848 14055 4868
rect 13759 3836 14055 3856
rect 13815 3834 13839 3836
rect 13895 3834 13919 3836
rect 13975 3834 13999 3836
rect 13837 3782 13839 3834
rect 13901 3782 13913 3834
rect 13975 3782 13977 3834
rect 13815 3780 13839 3782
rect 13895 3780 13919 3782
rect 13975 3780 13999 3782
rect 13759 3760 14055 3780
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13556 3182 13676 3210
rect 13556 3126 13584 3182
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13544 3120 13596 3126
rect 13544 3062 13596 3068
rect 13464 2854 13492 3062
rect 13832 2990 13860 3334
rect 13924 3126 13952 3334
rect 14108 3126 14136 5510
rect 14200 5030 14228 9930
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14476 9518 14504 9862
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14292 6730 14320 8434
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14384 7342 14412 7822
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14384 6866 14412 7278
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14292 6338 14320 6666
rect 14476 6390 14504 9318
rect 14568 9178 14596 14214
rect 14660 12458 14688 15302
rect 14752 13977 14780 15914
rect 15212 15706 15240 16050
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14936 15162 14964 15438
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14844 14618 14872 14894
rect 15028 14890 15056 14962
rect 15016 14884 15068 14890
rect 15016 14826 15068 14832
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14738 13968 14794 13977
rect 14738 13903 14794 13912
rect 14832 13456 14884 13462
rect 14832 13398 14884 13404
rect 14660 12430 14780 12458
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 14660 12102 14688 12242
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 9994 14688 12038
rect 14648 9988 14700 9994
rect 14648 9930 14700 9936
rect 14752 9874 14780 12430
rect 14660 9846 14780 9874
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14660 7970 14688 9846
rect 14844 9738 14872 13398
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14936 12442 14964 13194
rect 15028 12986 15056 14826
rect 15304 14618 15332 16118
rect 15488 15638 15516 16546
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15672 16046 15700 16390
rect 15568 16040 15620 16046
rect 15568 15982 15620 15988
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15304 13938 15332 14554
rect 15580 14074 15608 15982
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15672 13938 15700 14350
rect 15752 14340 15804 14346
rect 15752 14282 15804 14288
rect 15764 13938 15792 14282
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 15120 12850 15148 13194
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15212 12730 15240 13126
rect 15488 12850 15516 13126
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15120 12702 15240 12730
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14936 11558 14964 11698
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14936 10674 14964 11494
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14936 10130 14964 10610
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14752 9710 14872 9738
rect 14752 9654 14780 9710
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 8974 14780 9454
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14660 7942 14780 7970
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14556 7404 14608 7410
rect 14660 7392 14688 7822
rect 14752 7546 14780 7942
rect 14844 7818 14872 9522
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 14832 7812 14884 7818
rect 14832 7754 14884 7760
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14608 7364 14688 7392
rect 14740 7404 14792 7410
rect 14556 7346 14608 7352
rect 14740 7346 14792 7352
rect 14568 7206 14596 7346
rect 14752 7290 14780 7346
rect 14660 7262 14780 7290
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14464 6384 14516 6390
rect 14292 6310 14412 6338
rect 14464 6326 14516 6332
rect 14280 6180 14332 6186
rect 14280 6122 14332 6128
rect 14292 5545 14320 6122
rect 14384 5710 14412 6310
rect 14568 5710 14596 7142
rect 14660 6458 14688 7262
rect 14648 6452 14700 6458
rect 14936 6440 14964 8842
rect 15028 6662 15056 12582
rect 15120 11830 15148 12702
rect 15488 12238 15516 12786
rect 15580 12238 15608 12786
rect 15672 12442 15700 13874
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15764 11898 15792 13874
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15108 11824 15160 11830
rect 15108 11766 15160 11772
rect 15120 10674 15148 11766
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15212 10538 15240 11494
rect 15764 11150 15792 11834
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15488 10810 15516 11086
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15120 8022 15148 9998
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15212 8498 15240 9522
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15212 8090 15240 8434
rect 15304 8430 15332 9522
rect 15660 8900 15712 8906
rect 15660 8842 15712 8848
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15672 8265 15700 8842
rect 15658 8256 15714 8265
rect 15658 8191 15714 8200
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15120 7410 15148 7958
rect 15292 7812 15344 7818
rect 15292 7754 15344 7760
rect 15304 7546 15332 7754
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14648 6394 14700 6400
rect 14844 6412 14964 6440
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14278 5536 14334 5545
rect 14278 5471 14334 5480
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4826 14228 4966
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14384 4622 14412 5646
rect 14568 5166 14596 5646
rect 14660 5642 14688 6394
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14372 4616 14424 4622
rect 14292 4576 14372 4604
rect 14292 4146 14320 4576
rect 14372 4558 14424 4564
rect 14568 4214 14596 5102
rect 14660 4622 14688 5578
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14752 4554 14780 5782
rect 14844 5778 14872 6412
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 14832 5772 14884 5778
rect 14832 5714 14884 5720
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14556 4208 14608 4214
rect 14556 4150 14608 4156
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14200 3602 14228 3878
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14292 3534 14320 3674
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13759 2748 14055 2768
rect 13815 2746 13839 2748
rect 13895 2746 13919 2748
rect 13975 2746 13999 2748
rect 13837 2694 13839 2746
rect 13901 2694 13913 2746
rect 13975 2694 13977 2746
rect 13815 2692 13839 2694
rect 13895 2692 13919 2694
rect 13975 2692 13999 2694
rect 13759 2672 14055 2692
rect 14384 2446 14412 4150
rect 14464 4004 14516 4010
rect 14464 3946 14516 3952
rect 14476 3466 14504 3946
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14752 2774 14780 4490
rect 14844 4078 14872 5714
rect 14936 5370 14964 6258
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 14936 4214 14964 5306
rect 15028 4690 15056 5714
rect 15120 5710 15148 7346
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15304 6254 15332 6734
rect 15396 6322 15424 6802
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 15028 4486 15056 4626
rect 15016 4480 15068 4486
rect 15016 4422 15068 4428
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14844 3754 14872 4014
rect 14844 3726 14964 3754
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14844 3126 14872 3538
rect 14936 3398 14964 3726
rect 15120 3534 15148 5170
rect 15212 4214 15240 5510
rect 15304 4282 15332 6190
rect 15384 5636 15436 5642
rect 15384 5578 15436 5584
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15200 4208 15252 4214
rect 15200 4150 15252 4156
rect 15396 3738 15424 5578
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14832 3120 14884 3126
rect 14832 3062 14884 3068
rect 15396 3058 15424 3674
rect 17500 3188 17552 3194
rect 17500 3130 17552 3136
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 14660 2746 14780 2774
rect 14660 2650 14688 2746
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 15764 2553 15792 2858
rect 15750 2544 15806 2553
rect 15750 2479 15806 2488
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 13360 2372 13412 2378
rect 13360 2314 13412 2320
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15660 2372 15712 2378
rect 15660 2314 15712 2320
rect 13372 870 13492 898
rect 13372 762 13400 870
rect 13464 800 13492 870
rect 15488 800 15516 2314
rect 15672 2038 15700 2314
rect 15660 2032 15712 2038
rect 15660 1974 15712 1980
rect 17512 800 17540 3130
rect 13004 734 13400 762
rect 13450 0 13506 800
rect 15474 0 15530 800
rect 17498 0 17554 800
<< via2 >>
rect 1858 17212 1860 17232
rect 1860 17212 1912 17232
rect 1912 17212 1914 17232
rect 1858 17176 1914 17212
rect 6077 17434 6133 17436
rect 6157 17434 6213 17436
rect 6237 17434 6293 17436
rect 6317 17434 6373 17436
rect 6077 17382 6103 17434
rect 6103 17382 6133 17434
rect 6157 17382 6167 17434
rect 6167 17382 6213 17434
rect 6237 17382 6283 17434
rect 6283 17382 6293 17434
rect 6317 17382 6347 17434
rect 6347 17382 6373 17434
rect 6077 17380 6133 17382
rect 6157 17380 6213 17382
rect 6237 17380 6293 17382
rect 6317 17380 6373 17382
rect 11198 17434 11254 17436
rect 11278 17434 11334 17436
rect 11358 17434 11414 17436
rect 11438 17434 11494 17436
rect 11198 17382 11224 17434
rect 11224 17382 11254 17434
rect 11278 17382 11288 17434
rect 11288 17382 11334 17434
rect 11358 17382 11404 17434
rect 11404 17382 11414 17434
rect 11438 17382 11468 17434
rect 11468 17382 11494 17434
rect 11198 17380 11254 17382
rect 11278 17380 11334 17382
rect 11358 17380 11414 17382
rect 11438 17380 11494 17382
rect 3516 16890 3572 16892
rect 3596 16890 3652 16892
rect 3676 16890 3732 16892
rect 3756 16890 3812 16892
rect 3516 16838 3542 16890
rect 3542 16838 3572 16890
rect 3596 16838 3606 16890
rect 3606 16838 3652 16890
rect 3676 16838 3722 16890
rect 3722 16838 3732 16890
rect 3756 16838 3786 16890
rect 3786 16838 3812 16890
rect 3516 16836 3572 16838
rect 3596 16836 3652 16838
rect 3676 16836 3732 16838
rect 3756 16836 3812 16838
rect 1950 14184 2006 14240
rect 1858 11464 1914 11520
rect 1398 5752 1454 5808
rect 1582 3032 1638 3088
rect 3516 15802 3572 15804
rect 3596 15802 3652 15804
rect 3676 15802 3732 15804
rect 3756 15802 3812 15804
rect 3516 15750 3542 15802
rect 3542 15750 3572 15802
rect 3596 15750 3606 15802
rect 3606 15750 3652 15802
rect 3676 15750 3722 15802
rect 3722 15750 3732 15802
rect 3756 15750 3786 15802
rect 3786 15750 3812 15802
rect 3516 15748 3572 15750
rect 3596 15748 3652 15750
rect 3676 15748 3732 15750
rect 3756 15748 3812 15750
rect 3516 14714 3572 14716
rect 3596 14714 3652 14716
rect 3676 14714 3732 14716
rect 3756 14714 3812 14716
rect 3516 14662 3542 14714
rect 3542 14662 3572 14714
rect 3596 14662 3606 14714
rect 3606 14662 3652 14714
rect 3676 14662 3722 14714
rect 3722 14662 3732 14714
rect 3756 14662 3786 14714
rect 3786 14662 3812 14714
rect 3516 14660 3572 14662
rect 3596 14660 3652 14662
rect 3676 14660 3732 14662
rect 3756 14660 3812 14662
rect 3516 13626 3572 13628
rect 3596 13626 3652 13628
rect 3676 13626 3732 13628
rect 3756 13626 3812 13628
rect 3516 13574 3542 13626
rect 3542 13574 3572 13626
rect 3596 13574 3606 13626
rect 3606 13574 3652 13626
rect 3676 13574 3722 13626
rect 3722 13574 3732 13626
rect 3756 13574 3786 13626
rect 3786 13574 3812 13626
rect 3516 13572 3572 13574
rect 3596 13572 3652 13574
rect 3676 13572 3732 13574
rect 3756 13572 3812 13574
rect 3516 12538 3572 12540
rect 3596 12538 3652 12540
rect 3676 12538 3732 12540
rect 3756 12538 3812 12540
rect 3516 12486 3542 12538
rect 3542 12486 3572 12538
rect 3596 12486 3606 12538
rect 3606 12486 3652 12538
rect 3676 12486 3722 12538
rect 3722 12486 3732 12538
rect 3756 12486 3786 12538
rect 3786 12486 3812 12538
rect 3516 12484 3572 12486
rect 3596 12484 3652 12486
rect 3676 12484 3732 12486
rect 3756 12484 3812 12486
rect 3516 11450 3572 11452
rect 3596 11450 3652 11452
rect 3676 11450 3732 11452
rect 3756 11450 3812 11452
rect 3516 11398 3542 11450
rect 3542 11398 3572 11450
rect 3596 11398 3606 11450
rect 3606 11398 3652 11450
rect 3676 11398 3722 11450
rect 3722 11398 3732 11450
rect 3756 11398 3786 11450
rect 3786 11398 3812 11450
rect 3516 11396 3572 11398
rect 3596 11396 3652 11398
rect 3676 11396 3732 11398
rect 3756 11396 3812 11398
rect 3516 10362 3572 10364
rect 3596 10362 3652 10364
rect 3676 10362 3732 10364
rect 3756 10362 3812 10364
rect 3516 10310 3542 10362
rect 3542 10310 3572 10362
rect 3596 10310 3606 10362
rect 3606 10310 3652 10362
rect 3676 10310 3722 10362
rect 3722 10310 3732 10362
rect 3756 10310 3786 10362
rect 3786 10310 3812 10362
rect 3516 10308 3572 10310
rect 3596 10308 3652 10310
rect 3676 10308 3732 10310
rect 3756 10308 3812 10310
rect 3516 9274 3572 9276
rect 3596 9274 3652 9276
rect 3676 9274 3732 9276
rect 3756 9274 3812 9276
rect 3516 9222 3542 9274
rect 3542 9222 3572 9274
rect 3596 9222 3606 9274
rect 3606 9222 3652 9274
rect 3676 9222 3722 9274
rect 3722 9222 3732 9274
rect 3756 9222 3786 9274
rect 3786 9222 3812 9274
rect 3516 9220 3572 9222
rect 3596 9220 3652 9222
rect 3676 9220 3732 9222
rect 3756 9220 3812 9222
rect 2870 8472 2926 8528
rect 3516 8186 3572 8188
rect 3596 8186 3652 8188
rect 3676 8186 3732 8188
rect 3756 8186 3812 8188
rect 3516 8134 3542 8186
rect 3542 8134 3572 8186
rect 3596 8134 3606 8186
rect 3606 8134 3652 8186
rect 3676 8134 3722 8186
rect 3722 8134 3732 8186
rect 3756 8134 3786 8186
rect 3786 8134 3812 8186
rect 3516 8132 3572 8134
rect 3596 8132 3652 8134
rect 3676 8132 3732 8134
rect 3756 8132 3812 8134
rect 3516 7098 3572 7100
rect 3596 7098 3652 7100
rect 3676 7098 3732 7100
rect 3756 7098 3812 7100
rect 3516 7046 3542 7098
rect 3542 7046 3572 7098
rect 3596 7046 3606 7098
rect 3606 7046 3652 7098
rect 3676 7046 3722 7098
rect 3722 7046 3732 7098
rect 3756 7046 3786 7098
rect 3786 7046 3812 7098
rect 3516 7044 3572 7046
rect 3596 7044 3652 7046
rect 3676 7044 3732 7046
rect 3756 7044 3812 7046
rect 2502 5752 2558 5808
rect 2778 5752 2834 5808
rect 3516 6010 3572 6012
rect 3596 6010 3652 6012
rect 3676 6010 3732 6012
rect 3756 6010 3812 6012
rect 3516 5958 3542 6010
rect 3542 5958 3572 6010
rect 3596 5958 3606 6010
rect 3606 5958 3652 6010
rect 3676 5958 3722 6010
rect 3722 5958 3732 6010
rect 3756 5958 3786 6010
rect 3786 5958 3812 6010
rect 3516 5956 3572 5958
rect 3596 5956 3652 5958
rect 3676 5956 3732 5958
rect 3756 5956 3812 5958
rect 2686 3440 2742 3496
rect 2594 3188 2650 3224
rect 2594 3168 2596 3188
rect 2596 3168 2648 3188
rect 2648 3168 2650 3188
rect 2778 2760 2834 2816
rect 3516 4922 3572 4924
rect 3596 4922 3652 4924
rect 3676 4922 3732 4924
rect 3756 4922 3812 4924
rect 3516 4870 3542 4922
rect 3542 4870 3572 4922
rect 3596 4870 3606 4922
rect 3606 4870 3652 4922
rect 3676 4870 3722 4922
rect 3722 4870 3732 4922
rect 3756 4870 3786 4922
rect 3786 4870 3812 4922
rect 3516 4868 3572 4870
rect 3596 4868 3652 4870
rect 3676 4868 3732 4870
rect 3756 4868 3812 4870
rect 3516 3834 3572 3836
rect 3596 3834 3652 3836
rect 3676 3834 3732 3836
rect 3756 3834 3812 3836
rect 3516 3782 3542 3834
rect 3542 3782 3572 3834
rect 3596 3782 3606 3834
rect 3606 3782 3652 3834
rect 3676 3782 3722 3834
rect 3722 3782 3732 3834
rect 3756 3782 3786 3834
rect 3786 3782 3812 3834
rect 3516 3780 3572 3782
rect 3596 3780 3652 3782
rect 3676 3780 3732 3782
rect 3756 3780 3812 3782
rect 3882 3576 3938 3632
rect 6077 16346 6133 16348
rect 6157 16346 6213 16348
rect 6237 16346 6293 16348
rect 6317 16346 6373 16348
rect 6077 16294 6103 16346
rect 6103 16294 6133 16346
rect 6157 16294 6167 16346
rect 6167 16294 6213 16346
rect 6237 16294 6283 16346
rect 6283 16294 6293 16346
rect 6317 16294 6347 16346
rect 6347 16294 6373 16346
rect 6077 16292 6133 16294
rect 6157 16292 6213 16294
rect 6237 16292 6293 16294
rect 6317 16292 6373 16294
rect 6077 15258 6133 15260
rect 6157 15258 6213 15260
rect 6237 15258 6293 15260
rect 6317 15258 6373 15260
rect 6077 15206 6103 15258
rect 6103 15206 6133 15258
rect 6157 15206 6167 15258
rect 6167 15206 6213 15258
rect 6237 15206 6283 15258
rect 6283 15206 6293 15258
rect 6317 15206 6347 15258
rect 6347 15206 6373 15258
rect 6077 15204 6133 15206
rect 6157 15204 6213 15206
rect 6237 15204 6293 15206
rect 6317 15204 6373 15206
rect 6077 14170 6133 14172
rect 6157 14170 6213 14172
rect 6237 14170 6293 14172
rect 6317 14170 6373 14172
rect 6077 14118 6103 14170
rect 6103 14118 6133 14170
rect 6157 14118 6167 14170
rect 6167 14118 6213 14170
rect 6237 14118 6283 14170
rect 6283 14118 6293 14170
rect 6317 14118 6347 14170
rect 6347 14118 6373 14170
rect 6077 14116 6133 14118
rect 6157 14116 6213 14118
rect 6237 14116 6293 14118
rect 6317 14116 6373 14118
rect 6077 13082 6133 13084
rect 6157 13082 6213 13084
rect 6237 13082 6293 13084
rect 6317 13082 6373 13084
rect 6077 13030 6103 13082
rect 6103 13030 6133 13082
rect 6157 13030 6167 13082
rect 6167 13030 6213 13082
rect 6237 13030 6283 13082
rect 6283 13030 6293 13082
rect 6317 13030 6347 13082
rect 6347 13030 6373 13082
rect 6077 13028 6133 13030
rect 6157 13028 6213 13030
rect 6237 13028 6293 13030
rect 6317 13028 6373 13030
rect 8638 16890 8694 16892
rect 8718 16890 8774 16892
rect 8798 16890 8854 16892
rect 8878 16890 8934 16892
rect 8638 16838 8664 16890
rect 8664 16838 8694 16890
rect 8718 16838 8728 16890
rect 8728 16838 8774 16890
rect 8798 16838 8844 16890
rect 8844 16838 8854 16890
rect 8878 16838 8908 16890
rect 8908 16838 8934 16890
rect 8638 16836 8694 16838
rect 8718 16836 8774 16838
rect 8798 16836 8854 16838
rect 8878 16836 8934 16838
rect 5354 7928 5410 7984
rect 4618 7404 4674 7440
rect 4618 7384 4620 7404
rect 4620 7384 4672 7404
rect 4672 7384 4674 7404
rect 4802 7268 4858 7304
rect 4802 7248 4804 7268
rect 4804 7248 4856 7268
rect 4856 7248 4858 7268
rect 6077 11994 6133 11996
rect 6157 11994 6213 11996
rect 6237 11994 6293 11996
rect 6317 11994 6373 11996
rect 6077 11942 6103 11994
rect 6103 11942 6133 11994
rect 6157 11942 6167 11994
rect 6167 11942 6213 11994
rect 6237 11942 6283 11994
rect 6283 11942 6293 11994
rect 6317 11942 6347 11994
rect 6347 11942 6373 11994
rect 6077 11940 6133 11942
rect 6157 11940 6213 11942
rect 6237 11940 6293 11942
rect 6317 11940 6373 11942
rect 6077 10906 6133 10908
rect 6157 10906 6213 10908
rect 6237 10906 6293 10908
rect 6317 10906 6373 10908
rect 6077 10854 6103 10906
rect 6103 10854 6133 10906
rect 6157 10854 6167 10906
rect 6167 10854 6213 10906
rect 6237 10854 6283 10906
rect 6283 10854 6293 10906
rect 6317 10854 6347 10906
rect 6347 10854 6373 10906
rect 6077 10852 6133 10854
rect 6157 10852 6213 10854
rect 6237 10852 6293 10854
rect 6317 10852 6373 10854
rect 6077 9818 6133 9820
rect 6157 9818 6213 9820
rect 6237 9818 6293 9820
rect 6317 9818 6373 9820
rect 6077 9766 6103 9818
rect 6103 9766 6133 9818
rect 6157 9766 6167 9818
rect 6167 9766 6213 9818
rect 6237 9766 6283 9818
rect 6283 9766 6293 9818
rect 6317 9766 6347 9818
rect 6347 9766 6373 9818
rect 6077 9764 6133 9766
rect 6157 9764 6213 9766
rect 6237 9764 6293 9766
rect 6317 9764 6373 9766
rect 5354 6840 5410 6896
rect 4434 2932 4436 2952
rect 4436 2932 4488 2952
rect 4488 2932 4490 2952
rect 4434 2896 4490 2932
rect 3516 2746 3572 2748
rect 3596 2746 3652 2748
rect 3676 2746 3732 2748
rect 3756 2746 3812 2748
rect 3516 2694 3542 2746
rect 3542 2694 3572 2746
rect 3596 2694 3606 2746
rect 3606 2694 3652 2746
rect 3676 2694 3722 2746
rect 3722 2694 3732 2746
rect 3756 2694 3786 2746
rect 3786 2694 3812 2746
rect 3516 2692 3572 2694
rect 3596 2692 3652 2694
rect 3676 2692 3732 2694
rect 3756 2692 3812 2694
rect 5630 3168 5686 3224
rect 6077 8730 6133 8732
rect 6157 8730 6213 8732
rect 6237 8730 6293 8732
rect 6317 8730 6373 8732
rect 6077 8678 6103 8730
rect 6103 8678 6133 8730
rect 6157 8678 6167 8730
rect 6167 8678 6213 8730
rect 6237 8678 6283 8730
rect 6283 8678 6293 8730
rect 6317 8678 6347 8730
rect 6347 8678 6373 8730
rect 6077 8676 6133 8678
rect 6157 8676 6213 8678
rect 6237 8676 6293 8678
rect 6317 8676 6373 8678
rect 6077 7642 6133 7644
rect 6157 7642 6213 7644
rect 6237 7642 6293 7644
rect 6317 7642 6373 7644
rect 6077 7590 6103 7642
rect 6103 7590 6133 7642
rect 6157 7590 6167 7642
rect 6167 7590 6213 7642
rect 6237 7590 6283 7642
rect 6283 7590 6293 7642
rect 6317 7590 6347 7642
rect 6347 7590 6373 7642
rect 6077 7588 6133 7590
rect 6157 7588 6213 7590
rect 6237 7588 6293 7590
rect 6317 7588 6373 7590
rect 6077 6554 6133 6556
rect 6157 6554 6213 6556
rect 6237 6554 6293 6556
rect 6317 6554 6373 6556
rect 6077 6502 6103 6554
rect 6103 6502 6133 6554
rect 6157 6502 6167 6554
rect 6167 6502 6213 6554
rect 6237 6502 6283 6554
rect 6283 6502 6293 6554
rect 6317 6502 6347 6554
rect 6347 6502 6373 6554
rect 6077 6500 6133 6502
rect 6157 6500 6213 6502
rect 6237 6500 6293 6502
rect 6317 6500 6373 6502
rect 6550 7792 6606 7848
rect 6642 7656 6698 7712
rect 6642 6568 6698 6624
rect 6458 6296 6514 6352
rect 5906 5888 5962 5944
rect 6077 5466 6133 5468
rect 6157 5466 6213 5468
rect 6237 5466 6293 5468
rect 6317 5466 6373 5468
rect 6077 5414 6103 5466
rect 6103 5414 6133 5466
rect 6157 5414 6167 5466
rect 6167 5414 6213 5466
rect 6237 5414 6283 5466
rect 6283 5414 6293 5466
rect 6317 5414 6347 5466
rect 6347 5414 6373 5466
rect 6077 5412 6133 5414
rect 6157 5412 6213 5414
rect 6237 5412 6293 5414
rect 6317 5412 6373 5414
rect 7010 6976 7066 7032
rect 8638 15802 8694 15804
rect 8718 15802 8774 15804
rect 8798 15802 8854 15804
rect 8878 15802 8934 15804
rect 8638 15750 8664 15802
rect 8664 15750 8694 15802
rect 8718 15750 8728 15802
rect 8728 15750 8774 15802
rect 8798 15750 8844 15802
rect 8844 15750 8854 15802
rect 8878 15750 8908 15802
rect 8908 15750 8934 15802
rect 8638 15748 8694 15750
rect 8718 15748 8774 15750
rect 8798 15748 8854 15750
rect 8878 15748 8934 15750
rect 11198 16346 11254 16348
rect 11278 16346 11334 16348
rect 11358 16346 11414 16348
rect 11438 16346 11494 16348
rect 11198 16294 11224 16346
rect 11224 16294 11254 16346
rect 11278 16294 11288 16346
rect 11288 16294 11334 16346
rect 11358 16294 11404 16346
rect 11404 16294 11414 16346
rect 11438 16294 11468 16346
rect 11468 16294 11494 16346
rect 11198 16292 11254 16294
rect 11278 16292 11334 16294
rect 11358 16292 11414 16294
rect 11438 16292 11494 16294
rect 8638 14714 8694 14716
rect 8718 14714 8774 14716
rect 8798 14714 8854 14716
rect 8878 14714 8934 14716
rect 8638 14662 8664 14714
rect 8664 14662 8694 14714
rect 8718 14662 8728 14714
rect 8728 14662 8774 14714
rect 8798 14662 8844 14714
rect 8844 14662 8854 14714
rect 8878 14662 8908 14714
rect 8908 14662 8934 14714
rect 8638 14660 8694 14662
rect 8718 14660 8774 14662
rect 8798 14660 8854 14662
rect 8878 14660 8934 14662
rect 8638 13626 8694 13628
rect 8718 13626 8774 13628
rect 8798 13626 8854 13628
rect 8878 13626 8934 13628
rect 8638 13574 8664 13626
rect 8664 13574 8694 13626
rect 8718 13574 8728 13626
rect 8728 13574 8774 13626
rect 8798 13574 8844 13626
rect 8844 13574 8854 13626
rect 8878 13574 8908 13626
rect 8908 13574 8934 13626
rect 8638 13572 8694 13574
rect 8718 13572 8774 13574
rect 8798 13572 8854 13574
rect 8878 13572 8934 13574
rect 8638 12538 8694 12540
rect 8718 12538 8774 12540
rect 8798 12538 8854 12540
rect 8878 12538 8934 12540
rect 8638 12486 8664 12538
rect 8664 12486 8694 12538
rect 8718 12486 8728 12538
rect 8728 12486 8774 12538
rect 8798 12486 8844 12538
rect 8844 12486 8854 12538
rect 8878 12486 8908 12538
rect 8908 12486 8934 12538
rect 8638 12484 8694 12486
rect 8718 12484 8774 12486
rect 8798 12484 8854 12486
rect 8878 12484 8934 12486
rect 6077 4378 6133 4380
rect 6157 4378 6213 4380
rect 6237 4378 6293 4380
rect 6317 4378 6373 4380
rect 6077 4326 6103 4378
rect 6103 4326 6133 4378
rect 6157 4326 6167 4378
rect 6167 4326 6213 4378
rect 6237 4326 6283 4378
rect 6283 4326 6293 4378
rect 6317 4326 6347 4378
rect 6347 4326 6373 4378
rect 6077 4324 6133 4326
rect 6157 4324 6213 4326
rect 6237 4324 6293 4326
rect 6317 4324 6373 4326
rect 7286 4256 7342 4312
rect 6090 3476 6092 3496
rect 6092 3476 6144 3496
rect 6144 3476 6146 3496
rect 6090 3440 6146 3476
rect 6077 3290 6133 3292
rect 6157 3290 6213 3292
rect 6237 3290 6293 3292
rect 6317 3290 6373 3292
rect 6077 3238 6103 3290
rect 6103 3238 6133 3290
rect 6157 3238 6167 3290
rect 6167 3238 6213 3290
rect 6237 3238 6283 3290
rect 6283 3238 6293 3290
rect 6317 3238 6347 3290
rect 6347 3238 6373 3290
rect 6077 3236 6133 3238
rect 6157 3236 6213 3238
rect 6237 3236 6293 3238
rect 6317 3236 6373 3238
rect 7102 3984 7158 4040
rect 7194 3460 7250 3496
rect 7194 3440 7196 3460
rect 7196 3440 7248 3460
rect 7248 3440 7250 3460
rect 7102 3032 7158 3088
rect 7286 3068 7288 3088
rect 7288 3068 7340 3088
rect 7340 3068 7342 3088
rect 7286 3032 7342 3068
rect 7010 2916 7066 2952
rect 7010 2896 7012 2916
rect 7012 2896 7064 2916
rect 7064 2896 7066 2916
rect 6077 2202 6133 2204
rect 6157 2202 6213 2204
rect 6237 2202 6293 2204
rect 6317 2202 6373 2204
rect 6077 2150 6103 2202
rect 6103 2150 6133 2202
rect 6157 2150 6167 2202
rect 6167 2150 6213 2202
rect 6237 2150 6283 2202
rect 6283 2150 6293 2202
rect 6317 2150 6347 2202
rect 6347 2150 6373 2202
rect 6077 2148 6133 2150
rect 6157 2148 6213 2150
rect 6237 2148 6293 2150
rect 6317 2148 6373 2150
rect 7470 7540 7526 7576
rect 7470 7520 7472 7540
rect 7472 7520 7524 7540
rect 7524 7520 7526 7540
rect 7470 6740 7472 6760
rect 7472 6740 7524 6760
rect 7524 6740 7526 6760
rect 7470 6704 7526 6740
rect 7654 6604 7656 6624
rect 7656 6604 7708 6624
rect 7708 6604 7710 6624
rect 7654 6568 7710 6604
rect 8638 11450 8694 11452
rect 8718 11450 8774 11452
rect 8798 11450 8854 11452
rect 8878 11450 8934 11452
rect 8638 11398 8664 11450
rect 8664 11398 8694 11450
rect 8718 11398 8728 11450
rect 8728 11398 8774 11450
rect 8798 11398 8844 11450
rect 8844 11398 8854 11450
rect 8878 11398 8908 11450
rect 8908 11398 8934 11450
rect 8638 11396 8694 11398
rect 8718 11396 8774 11398
rect 8798 11396 8854 11398
rect 8878 11396 8934 11398
rect 11198 15258 11254 15260
rect 11278 15258 11334 15260
rect 11358 15258 11414 15260
rect 11438 15258 11494 15260
rect 11198 15206 11224 15258
rect 11224 15206 11254 15258
rect 11278 15206 11288 15258
rect 11288 15206 11334 15258
rect 11358 15206 11404 15258
rect 11404 15206 11414 15258
rect 11438 15206 11468 15258
rect 11468 15206 11494 15258
rect 11198 15204 11254 15206
rect 11278 15204 11334 15206
rect 11358 15204 11414 15206
rect 11438 15204 11494 15206
rect 11198 14170 11254 14172
rect 11278 14170 11334 14172
rect 11358 14170 11414 14172
rect 11438 14170 11494 14172
rect 11198 14118 11224 14170
rect 11224 14118 11254 14170
rect 11278 14118 11288 14170
rect 11288 14118 11334 14170
rect 11358 14118 11404 14170
rect 11404 14118 11414 14170
rect 11438 14118 11468 14170
rect 11468 14118 11494 14170
rect 11198 14116 11254 14118
rect 11278 14116 11334 14118
rect 11358 14116 11414 14118
rect 11438 14116 11494 14118
rect 8638 10362 8694 10364
rect 8718 10362 8774 10364
rect 8798 10362 8854 10364
rect 8878 10362 8934 10364
rect 8638 10310 8664 10362
rect 8664 10310 8694 10362
rect 8718 10310 8728 10362
rect 8728 10310 8774 10362
rect 8798 10310 8844 10362
rect 8844 10310 8854 10362
rect 8878 10310 8908 10362
rect 8908 10310 8934 10362
rect 8638 10308 8694 10310
rect 8718 10308 8774 10310
rect 8798 10308 8854 10310
rect 8878 10308 8934 10310
rect 8638 9274 8694 9276
rect 8718 9274 8774 9276
rect 8798 9274 8854 9276
rect 8878 9274 8934 9276
rect 8638 9222 8664 9274
rect 8664 9222 8694 9274
rect 8718 9222 8728 9274
rect 8728 9222 8774 9274
rect 8798 9222 8844 9274
rect 8844 9222 8854 9274
rect 8878 9222 8908 9274
rect 8908 9222 8934 9274
rect 8638 9220 8694 9222
rect 8718 9220 8774 9222
rect 8798 9220 8854 9222
rect 8878 9220 8934 9222
rect 8022 7112 8078 7168
rect 8638 8186 8694 8188
rect 8718 8186 8774 8188
rect 8798 8186 8854 8188
rect 8878 8186 8934 8188
rect 8638 8134 8664 8186
rect 8664 8134 8694 8186
rect 8718 8134 8728 8186
rect 8728 8134 8774 8186
rect 8798 8134 8844 8186
rect 8844 8134 8854 8186
rect 8878 8134 8908 8186
rect 8908 8134 8934 8186
rect 8638 8132 8694 8134
rect 8718 8132 8774 8134
rect 8798 8132 8854 8134
rect 8878 8132 8934 8134
rect 8390 7656 8446 7712
rect 8298 7520 8354 7576
rect 8482 7112 8538 7168
rect 8638 7098 8694 7100
rect 8718 7098 8774 7100
rect 8798 7098 8854 7100
rect 8878 7098 8934 7100
rect 8638 7046 8664 7098
rect 8664 7046 8694 7098
rect 8718 7046 8728 7098
rect 8728 7046 8774 7098
rect 8798 7046 8844 7098
rect 8844 7046 8854 7098
rect 8878 7046 8908 7098
rect 8908 7046 8934 7098
rect 8638 7044 8694 7046
rect 8718 7044 8774 7046
rect 8798 7044 8854 7046
rect 8878 7044 8934 7046
rect 8482 6976 8538 7032
rect 7930 6704 7986 6760
rect 7838 6432 7894 6488
rect 9126 6840 9182 6896
rect 8638 6010 8694 6012
rect 8718 6010 8774 6012
rect 8798 6010 8854 6012
rect 8878 6010 8934 6012
rect 8638 5958 8664 6010
rect 8664 5958 8694 6010
rect 8718 5958 8728 6010
rect 8728 5958 8774 6010
rect 8798 5958 8844 6010
rect 8844 5958 8854 6010
rect 8878 5958 8908 6010
rect 8908 5958 8934 6010
rect 8638 5956 8694 5958
rect 8718 5956 8774 5958
rect 8798 5956 8854 5958
rect 8878 5956 8934 5958
rect 8206 5888 8262 5944
rect 8390 4256 8446 4312
rect 7746 3576 7802 3632
rect 8206 4120 8262 4176
rect 8298 3984 8354 4040
rect 8298 3440 8354 3496
rect 8638 4922 8694 4924
rect 8718 4922 8774 4924
rect 8798 4922 8854 4924
rect 8878 4922 8934 4924
rect 8638 4870 8664 4922
rect 8664 4870 8694 4922
rect 8718 4870 8728 4922
rect 8728 4870 8774 4922
rect 8798 4870 8844 4922
rect 8844 4870 8854 4922
rect 8878 4870 8908 4922
rect 8908 4870 8934 4922
rect 8638 4868 8694 4870
rect 8718 4868 8774 4870
rect 8798 4868 8854 4870
rect 8878 4868 8934 4870
rect 9218 4256 9274 4312
rect 8638 3834 8694 3836
rect 8718 3834 8774 3836
rect 8798 3834 8854 3836
rect 8878 3834 8934 3836
rect 8638 3782 8664 3834
rect 8664 3782 8694 3834
rect 8718 3782 8728 3834
rect 8728 3782 8774 3834
rect 8798 3782 8844 3834
rect 8844 3782 8854 3834
rect 8878 3782 8908 3834
rect 8908 3782 8934 3834
rect 8638 3780 8694 3782
rect 8718 3780 8774 3782
rect 8798 3780 8854 3782
rect 8878 3780 8934 3782
rect 8758 3068 8760 3088
rect 8760 3068 8812 3088
rect 8812 3068 8814 3088
rect 8758 3032 8814 3068
rect 8638 2746 8694 2748
rect 8718 2746 8774 2748
rect 8798 2746 8854 2748
rect 8878 2746 8934 2748
rect 8638 2694 8664 2746
rect 8664 2694 8694 2746
rect 8718 2694 8728 2746
rect 8728 2694 8774 2746
rect 8798 2694 8844 2746
rect 8844 2694 8854 2746
rect 8878 2694 8908 2746
rect 8908 2694 8934 2746
rect 8638 2692 8694 2694
rect 8718 2692 8774 2694
rect 8798 2692 8854 2694
rect 8878 2692 8934 2694
rect 9402 4140 9458 4176
rect 9402 4120 9404 4140
rect 9404 4120 9456 4140
rect 9456 4120 9458 4140
rect 9862 7792 9918 7848
rect 9678 6704 9734 6760
rect 9770 6432 9826 6488
rect 9770 6180 9826 6216
rect 9770 6160 9772 6180
rect 9772 6160 9824 6180
rect 9824 6160 9826 6180
rect 10138 6432 10194 6488
rect 10322 6432 10378 6488
rect 10322 6296 10378 6352
rect 11198 13082 11254 13084
rect 11278 13082 11334 13084
rect 11358 13082 11414 13084
rect 11438 13082 11494 13084
rect 11198 13030 11224 13082
rect 11224 13030 11254 13082
rect 11278 13030 11288 13082
rect 11288 13030 11334 13082
rect 11358 13030 11404 13082
rect 11404 13030 11414 13082
rect 11438 13030 11468 13082
rect 11468 13030 11494 13082
rect 11198 13028 11254 13030
rect 11278 13028 11334 13030
rect 11358 13028 11414 13030
rect 11438 13028 11494 13030
rect 11198 11994 11254 11996
rect 11278 11994 11334 11996
rect 11358 11994 11414 11996
rect 11438 11994 11494 11996
rect 11198 11942 11224 11994
rect 11224 11942 11254 11994
rect 11278 11942 11288 11994
rect 11288 11942 11334 11994
rect 11358 11942 11404 11994
rect 11404 11942 11414 11994
rect 11438 11942 11468 11994
rect 11468 11942 11494 11994
rect 11198 11940 11254 11942
rect 11278 11940 11334 11942
rect 11358 11940 11414 11942
rect 11438 11940 11494 11942
rect 11198 10906 11254 10908
rect 11278 10906 11334 10908
rect 11358 10906 11414 10908
rect 11438 10906 11494 10908
rect 11198 10854 11224 10906
rect 11224 10854 11254 10906
rect 11278 10854 11288 10906
rect 11288 10854 11334 10906
rect 11358 10854 11404 10906
rect 11404 10854 11414 10906
rect 11438 10854 11468 10906
rect 11468 10854 11494 10906
rect 11198 10852 11254 10854
rect 11278 10852 11334 10854
rect 11358 10852 11414 10854
rect 11438 10852 11494 10854
rect 11198 9818 11254 9820
rect 11278 9818 11334 9820
rect 11358 9818 11414 9820
rect 11438 9818 11494 9820
rect 11198 9766 11224 9818
rect 11224 9766 11254 9818
rect 11278 9766 11288 9818
rect 11288 9766 11334 9818
rect 11358 9766 11404 9818
rect 11404 9766 11414 9818
rect 11438 9766 11468 9818
rect 11468 9766 11494 9818
rect 11198 9764 11254 9766
rect 11278 9764 11334 9766
rect 11358 9764 11414 9766
rect 11438 9764 11494 9766
rect 11198 8730 11254 8732
rect 11278 8730 11334 8732
rect 11358 8730 11414 8732
rect 11438 8730 11494 8732
rect 11198 8678 11224 8730
rect 11224 8678 11254 8730
rect 11278 8678 11288 8730
rect 11288 8678 11334 8730
rect 11358 8678 11404 8730
rect 11404 8678 11414 8730
rect 11438 8678 11468 8730
rect 11468 8678 11494 8730
rect 11198 8676 11254 8678
rect 11278 8676 11334 8678
rect 11358 8676 11414 8678
rect 11438 8676 11494 8678
rect 11198 7642 11254 7644
rect 11278 7642 11334 7644
rect 11358 7642 11414 7644
rect 11438 7642 11494 7644
rect 11198 7590 11224 7642
rect 11224 7590 11254 7642
rect 11278 7590 11288 7642
rect 11288 7590 11334 7642
rect 11358 7590 11404 7642
rect 11404 7590 11414 7642
rect 11438 7590 11468 7642
rect 11468 7590 11494 7642
rect 11198 7588 11254 7590
rect 11278 7588 11334 7590
rect 11358 7588 11414 7590
rect 11438 7588 11494 7590
rect 11150 7384 11206 7440
rect 10966 6976 11022 7032
rect 11518 7248 11574 7304
rect 11426 6840 11482 6896
rect 11198 6554 11254 6556
rect 11278 6554 11334 6556
rect 11358 6554 11414 6556
rect 11438 6554 11494 6556
rect 11198 6502 11224 6554
rect 11224 6502 11254 6554
rect 11278 6502 11288 6554
rect 11288 6502 11334 6554
rect 11358 6502 11404 6554
rect 11404 6502 11414 6554
rect 11438 6502 11468 6554
rect 11468 6502 11494 6554
rect 11198 6500 11254 6502
rect 11278 6500 11334 6502
rect 11358 6500 11414 6502
rect 11438 6500 11494 6502
rect 11198 5466 11254 5468
rect 11278 5466 11334 5468
rect 11358 5466 11414 5468
rect 11438 5466 11494 5468
rect 11198 5414 11224 5466
rect 11224 5414 11254 5466
rect 11278 5414 11288 5466
rect 11288 5414 11334 5466
rect 11358 5414 11404 5466
rect 11404 5414 11414 5466
rect 11438 5414 11468 5466
rect 11468 5414 11494 5466
rect 11198 5412 11254 5414
rect 11278 5412 11334 5414
rect 11358 5412 11414 5414
rect 11438 5412 11494 5414
rect 11794 6740 11796 6760
rect 11796 6740 11848 6760
rect 11848 6740 11850 6760
rect 11794 6704 11850 6740
rect 11794 6296 11850 6352
rect 11198 4378 11254 4380
rect 11278 4378 11334 4380
rect 11358 4378 11414 4380
rect 11438 4378 11494 4380
rect 11198 4326 11224 4378
rect 11224 4326 11254 4378
rect 11278 4326 11288 4378
rect 11288 4326 11334 4378
rect 11358 4326 11404 4378
rect 11404 4326 11414 4378
rect 11438 4326 11468 4378
rect 11468 4326 11494 4378
rect 11198 4324 11254 4326
rect 11278 4324 11334 4326
rect 11358 4324 11414 4326
rect 11438 4324 11494 4326
rect 11198 3290 11254 3292
rect 11278 3290 11334 3292
rect 11358 3290 11414 3292
rect 11438 3290 11494 3292
rect 11198 3238 11224 3290
rect 11224 3238 11254 3290
rect 11278 3238 11288 3290
rect 11288 3238 11334 3290
rect 11358 3238 11404 3290
rect 11404 3238 11414 3290
rect 11438 3238 11468 3290
rect 11468 3238 11494 3290
rect 11198 3236 11254 3238
rect 11278 3236 11334 3238
rect 11358 3236 11414 3238
rect 11438 3236 11494 3238
rect 10046 2896 10102 2952
rect 11198 2202 11254 2204
rect 11278 2202 11334 2204
rect 11358 2202 11414 2204
rect 11438 2202 11494 2204
rect 11198 2150 11224 2202
rect 11224 2150 11254 2202
rect 11278 2150 11288 2202
rect 11288 2150 11334 2202
rect 11358 2150 11404 2202
rect 11404 2150 11414 2202
rect 11438 2150 11468 2202
rect 11468 2150 11494 2202
rect 11198 2148 11254 2150
rect 11278 2148 11334 2150
rect 11358 2148 11414 2150
rect 11438 2148 11494 2150
rect 13759 16890 13815 16892
rect 13839 16890 13895 16892
rect 13919 16890 13975 16892
rect 13999 16890 14055 16892
rect 13759 16838 13785 16890
rect 13785 16838 13815 16890
rect 13839 16838 13849 16890
rect 13849 16838 13895 16890
rect 13919 16838 13965 16890
rect 13965 16838 13975 16890
rect 13999 16838 14029 16890
rect 14029 16838 14055 16890
rect 13759 16836 13815 16838
rect 13839 16836 13895 16838
rect 13919 16836 13975 16838
rect 13999 16836 14055 16838
rect 12530 11192 12586 11248
rect 12714 6976 12770 7032
rect 12990 7928 13046 7984
rect 12898 6840 12954 6896
rect 13759 15802 13815 15804
rect 13839 15802 13895 15804
rect 13919 15802 13975 15804
rect 13999 15802 14055 15804
rect 13759 15750 13785 15802
rect 13785 15750 13815 15802
rect 13839 15750 13849 15802
rect 13849 15750 13895 15802
rect 13919 15750 13965 15802
rect 13965 15750 13975 15802
rect 13999 15750 14029 15802
rect 14029 15750 14055 15802
rect 13759 15748 13815 15750
rect 13839 15748 13895 15750
rect 13919 15748 13975 15750
rect 13999 15748 14055 15750
rect 13759 14714 13815 14716
rect 13839 14714 13895 14716
rect 13919 14714 13975 14716
rect 13999 14714 14055 14716
rect 13759 14662 13785 14714
rect 13785 14662 13815 14714
rect 13839 14662 13849 14714
rect 13849 14662 13895 14714
rect 13919 14662 13965 14714
rect 13965 14662 13975 14714
rect 13999 14662 14029 14714
rect 14029 14662 14055 14714
rect 13759 14660 13815 14662
rect 13839 14660 13895 14662
rect 13919 14660 13975 14662
rect 13999 14660 14055 14662
rect 13759 13626 13815 13628
rect 13839 13626 13895 13628
rect 13919 13626 13975 13628
rect 13999 13626 14055 13628
rect 13759 13574 13785 13626
rect 13785 13574 13815 13626
rect 13839 13574 13849 13626
rect 13849 13574 13895 13626
rect 13919 13574 13965 13626
rect 13965 13574 13975 13626
rect 13999 13574 14029 13626
rect 14029 13574 14055 13626
rect 13759 13572 13815 13574
rect 13839 13572 13895 13574
rect 13919 13572 13975 13574
rect 13999 13572 14055 13574
rect 15750 16904 15806 16960
rect 13759 12538 13815 12540
rect 13839 12538 13895 12540
rect 13919 12538 13975 12540
rect 13999 12538 14055 12540
rect 13759 12486 13785 12538
rect 13785 12486 13815 12538
rect 13839 12486 13849 12538
rect 13849 12486 13895 12538
rect 13919 12486 13965 12538
rect 13965 12486 13975 12538
rect 13999 12486 14029 12538
rect 14029 12486 14055 12538
rect 13759 12484 13815 12486
rect 13839 12484 13895 12486
rect 13919 12484 13975 12486
rect 13999 12484 14055 12486
rect 13759 11450 13815 11452
rect 13839 11450 13895 11452
rect 13919 11450 13975 11452
rect 13999 11450 14055 11452
rect 13759 11398 13785 11450
rect 13785 11398 13815 11450
rect 13839 11398 13849 11450
rect 13849 11398 13895 11450
rect 13919 11398 13965 11450
rect 13965 11398 13975 11450
rect 13999 11398 14029 11450
rect 14029 11398 14055 11450
rect 13759 11396 13815 11398
rect 13839 11396 13895 11398
rect 13919 11396 13975 11398
rect 13999 11396 14055 11398
rect 13759 10362 13815 10364
rect 13839 10362 13895 10364
rect 13919 10362 13975 10364
rect 13999 10362 14055 10364
rect 13759 10310 13785 10362
rect 13785 10310 13815 10362
rect 13839 10310 13849 10362
rect 13849 10310 13895 10362
rect 13919 10310 13965 10362
rect 13965 10310 13975 10362
rect 13999 10310 14029 10362
rect 14029 10310 14055 10362
rect 13759 10308 13815 10310
rect 13839 10308 13895 10310
rect 13919 10308 13975 10310
rect 13999 10308 14055 10310
rect 13759 9274 13815 9276
rect 13839 9274 13895 9276
rect 13919 9274 13975 9276
rect 13999 9274 14055 9276
rect 13759 9222 13785 9274
rect 13785 9222 13815 9274
rect 13839 9222 13849 9274
rect 13849 9222 13895 9274
rect 13919 9222 13965 9274
rect 13965 9222 13975 9274
rect 13999 9222 14029 9274
rect 14029 9222 14055 9274
rect 13759 9220 13815 9222
rect 13839 9220 13895 9222
rect 13919 9220 13975 9222
rect 13999 9220 14055 9222
rect 13759 8186 13815 8188
rect 13839 8186 13895 8188
rect 13919 8186 13975 8188
rect 13999 8186 14055 8188
rect 13759 8134 13785 8186
rect 13785 8134 13815 8186
rect 13839 8134 13849 8186
rect 13849 8134 13895 8186
rect 13919 8134 13965 8186
rect 13965 8134 13975 8186
rect 13999 8134 14029 8186
rect 14029 8134 14055 8186
rect 13759 8132 13815 8134
rect 13839 8132 13895 8134
rect 13919 8132 13975 8134
rect 13999 8132 14055 8134
rect 13759 7098 13815 7100
rect 13839 7098 13895 7100
rect 13919 7098 13975 7100
rect 13999 7098 14055 7100
rect 13759 7046 13785 7098
rect 13785 7046 13815 7098
rect 13839 7046 13849 7098
rect 13849 7046 13895 7098
rect 13919 7046 13965 7098
rect 13965 7046 13975 7098
rect 13999 7046 14029 7098
rect 14029 7046 14055 7098
rect 13759 7044 13815 7046
rect 13839 7044 13895 7046
rect 13919 7044 13975 7046
rect 13999 7044 14055 7046
rect 13726 6160 13782 6216
rect 13759 6010 13815 6012
rect 13839 6010 13895 6012
rect 13919 6010 13975 6012
rect 13999 6010 14055 6012
rect 13759 5958 13785 6010
rect 13785 5958 13815 6010
rect 13839 5958 13849 6010
rect 13849 5958 13895 6010
rect 13919 5958 13965 6010
rect 13965 5958 13975 6010
rect 13999 5958 14029 6010
rect 14029 5958 14055 6010
rect 13759 5956 13815 5958
rect 13839 5956 13895 5958
rect 13919 5956 13975 5958
rect 13999 5956 14055 5958
rect 13759 4922 13815 4924
rect 13839 4922 13895 4924
rect 13919 4922 13975 4924
rect 13999 4922 14055 4924
rect 13759 4870 13785 4922
rect 13785 4870 13815 4922
rect 13839 4870 13849 4922
rect 13849 4870 13895 4922
rect 13919 4870 13965 4922
rect 13965 4870 13975 4922
rect 13999 4870 14029 4922
rect 14029 4870 14055 4922
rect 13759 4868 13815 4870
rect 13839 4868 13895 4870
rect 13919 4868 13975 4870
rect 13999 4868 14055 4870
rect 13759 3834 13815 3836
rect 13839 3834 13895 3836
rect 13919 3834 13975 3836
rect 13999 3834 14055 3836
rect 13759 3782 13785 3834
rect 13785 3782 13815 3834
rect 13839 3782 13849 3834
rect 13849 3782 13895 3834
rect 13919 3782 13965 3834
rect 13965 3782 13975 3834
rect 13999 3782 14029 3834
rect 14029 3782 14055 3834
rect 13759 3780 13815 3782
rect 13839 3780 13895 3782
rect 13919 3780 13975 3782
rect 13999 3780 14055 3782
rect 14738 13912 14794 13968
rect 15658 8200 15714 8256
rect 14278 5480 14334 5536
rect 13759 2746 13815 2748
rect 13839 2746 13895 2748
rect 13919 2746 13975 2748
rect 13999 2746 14055 2748
rect 13759 2694 13785 2746
rect 13785 2694 13815 2746
rect 13839 2694 13849 2746
rect 13849 2694 13895 2746
rect 13919 2694 13965 2746
rect 13965 2694 13975 2746
rect 13999 2694 14029 2746
rect 14029 2694 14055 2746
rect 13759 2692 13815 2694
rect 13839 2692 13895 2694
rect 13919 2692 13975 2694
rect 13999 2692 14055 2694
rect 15750 2488 15806 2544
<< metal3 >>
rect 6065 17440 6385 17441
rect 6065 17376 6073 17440
rect 6137 17376 6153 17440
rect 6217 17376 6233 17440
rect 6297 17376 6313 17440
rect 6377 17376 6385 17440
rect 6065 17375 6385 17376
rect 11186 17440 11506 17441
rect 11186 17376 11194 17440
rect 11258 17376 11274 17440
rect 11338 17376 11354 17440
rect 11418 17376 11434 17440
rect 11498 17376 11506 17440
rect 11186 17375 11506 17376
rect 0 17234 800 17264
rect 1853 17234 1919 17237
rect 0 17232 1919 17234
rect 0 17176 1858 17232
rect 1914 17176 1919 17232
rect 0 17174 1919 17176
rect 0 17144 800 17174
rect 1853 17171 1919 17174
rect 15745 16962 15811 16965
rect 16784 16962 17584 16992
rect 15745 16960 17584 16962
rect 15745 16904 15750 16960
rect 15806 16904 17584 16960
rect 15745 16902 17584 16904
rect 15745 16899 15811 16902
rect 3504 16896 3824 16897
rect 3504 16832 3512 16896
rect 3576 16832 3592 16896
rect 3656 16832 3672 16896
rect 3736 16832 3752 16896
rect 3816 16832 3824 16896
rect 3504 16831 3824 16832
rect 8626 16896 8946 16897
rect 8626 16832 8634 16896
rect 8698 16832 8714 16896
rect 8778 16832 8794 16896
rect 8858 16832 8874 16896
rect 8938 16832 8946 16896
rect 8626 16831 8946 16832
rect 13747 16896 14067 16897
rect 13747 16832 13755 16896
rect 13819 16832 13835 16896
rect 13899 16832 13915 16896
rect 13979 16832 13995 16896
rect 14059 16832 14067 16896
rect 16784 16872 17584 16902
rect 13747 16831 14067 16832
rect 6065 16352 6385 16353
rect 6065 16288 6073 16352
rect 6137 16288 6153 16352
rect 6217 16288 6233 16352
rect 6297 16288 6313 16352
rect 6377 16288 6385 16352
rect 6065 16287 6385 16288
rect 11186 16352 11506 16353
rect 11186 16288 11194 16352
rect 11258 16288 11274 16352
rect 11338 16288 11354 16352
rect 11418 16288 11434 16352
rect 11498 16288 11506 16352
rect 11186 16287 11506 16288
rect 3504 15808 3824 15809
rect 3504 15744 3512 15808
rect 3576 15744 3592 15808
rect 3656 15744 3672 15808
rect 3736 15744 3752 15808
rect 3816 15744 3824 15808
rect 3504 15743 3824 15744
rect 8626 15808 8946 15809
rect 8626 15744 8634 15808
rect 8698 15744 8714 15808
rect 8778 15744 8794 15808
rect 8858 15744 8874 15808
rect 8938 15744 8946 15808
rect 8626 15743 8946 15744
rect 13747 15808 14067 15809
rect 13747 15744 13755 15808
rect 13819 15744 13835 15808
rect 13899 15744 13915 15808
rect 13979 15744 13995 15808
rect 14059 15744 14067 15808
rect 13747 15743 14067 15744
rect 6065 15264 6385 15265
rect 6065 15200 6073 15264
rect 6137 15200 6153 15264
rect 6217 15200 6233 15264
rect 6297 15200 6313 15264
rect 6377 15200 6385 15264
rect 6065 15199 6385 15200
rect 11186 15264 11506 15265
rect 11186 15200 11194 15264
rect 11258 15200 11274 15264
rect 11338 15200 11354 15264
rect 11418 15200 11434 15264
rect 11498 15200 11506 15264
rect 11186 15199 11506 15200
rect 3504 14720 3824 14721
rect 3504 14656 3512 14720
rect 3576 14656 3592 14720
rect 3656 14656 3672 14720
rect 3736 14656 3752 14720
rect 3816 14656 3824 14720
rect 3504 14655 3824 14656
rect 8626 14720 8946 14721
rect 8626 14656 8634 14720
rect 8698 14656 8714 14720
rect 8778 14656 8794 14720
rect 8858 14656 8874 14720
rect 8938 14656 8946 14720
rect 8626 14655 8946 14656
rect 13747 14720 14067 14721
rect 13747 14656 13755 14720
rect 13819 14656 13835 14720
rect 13899 14656 13915 14720
rect 13979 14656 13995 14720
rect 14059 14656 14067 14720
rect 13747 14655 14067 14656
rect 0 14242 800 14272
rect 1945 14242 2011 14245
rect 0 14240 2011 14242
rect 0 14184 1950 14240
rect 2006 14184 2011 14240
rect 0 14182 2011 14184
rect 0 14152 800 14182
rect 1945 14179 2011 14182
rect 6065 14176 6385 14177
rect 6065 14112 6073 14176
rect 6137 14112 6153 14176
rect 6217 14112 6233 14176
rect 6297 14112 6313 14176
rect 6377 14112 6385 14176
rect 6065 14111 6385 14112
rect 11186 14176 11506 14177
rect 11186 14112 11194 14176
rect 11258 14112 11274 14176
rect 11338 14112 11354 14176
rect 11418 14112 11434 14176
rect 11498 14112 11506 14176
rect 11186 14111 11506 14112
rect 14733 13970 14799 13973
rect 16784 13970 17584 14000
rect 14733 13968 17584 13970
rect 14733 13912 14738 13968
rect 14794 13912 17584 13968
rect 14733 13910 17584 13912
rect 14733 13907 14799 13910
rect 16784 13880 17584 13910
rect 3504 13632 3824 13633
rect 3504 13568 3512 13632
rect 3576 13568 3592 13632
rect 3656 13568 3672 13632
rect 3736 13568 3752 13632
rect 3816 13568 3824 13632
rect 3504 13567 3824 13568
rect 8626 13632 8946 13633
rect 8626 13568 8634 13632
rect 8698 13568 8714 13632
rect 8778 13568 8794 13632
rect 8858 13568 8874 13632
rect 8938 13568 8946 13632
rect 8626 13567 8946 13568
rect 13747 13632 14067 13633
rect 13747 13568 13755 13632
rect 13819 13568 13835 13632
rect 13899 13568 13915 13632
rect 13979 13568 13995 13632
rect 14059 13568 14067 13632
rect 13747 13567 14067 13568
rect 6065 13088 6385 13089
rect 6065 13024 6073 13088
rect 6137 13024 6153 13088
rect 6217 13024 6233 13088
rect 6297 13024 6313 13088
rect 6377 13024 6385 13088
rect 6065 13023 6385 13024
rect 11186 13088 11506 13089
rect 11186 13024 11194 13088
rect 11258 13024 11274 13088
rect 11338 13024 11354 13088
rect 11418 13024 11434 13088
rect 11498 13024 11506 13088
rect 11186 13023 11506 13024
rect 3504 12544 3824 12545
rect 3504 12480 3512 12544
rect 3576 12480 3592 12544
rect 3656 12480 3672 12544
rect 3736 12480 3752 12544
rect 3816 12480 3824 12544
rect 3504 12479 3824 12480
rect 8626 12544 8946 12545
rect 8626 12480 8634 12544
rect 8698 12480 8714 12544
rect 8778 12480 8794 12544
rect 8858 12480 8874 12544
rect 8938 12480 8946 12544
rect 8626 12479 8946 12480
rect 13747 12544 14067 12545
rect 13747 12480 13755 12544
rect 13819 12480 13835 12544
rect 13899 12480 13915 12544
rect 13979 12480 13995 12544
rect 14059 12480 14067 12544
rect 13747 12479 14067 12480
rect 6065 12000 6385 12001
rect 6065 11936 6073 12000
rect 6137 11936 6153 12000
rect 6217 11936 6233 12000
rect 6297 11936 6313 12000
rect 6377 11936 6385 12000
rect 6065 11935 6385 11936
rect 11186 12000 11506 12001
rect 11186 11936 11194 12000
rect 11258 11936 11274 12000
rect 11338 11936 11354 12000
rect 11418 11936 11434 12000
rect 11498 11936 11506 12000
rect 11186 11935 11506 11936
rect 0 11522 800 11552
rect 1853 11522 1919 11525
rect 0 11520 1919 11522
rect 0 11464 1858 11520
rect 1914 11464 1919 11520
rect 0 11462 1919 11464
rect 0 11432 800 11462
rect 1853 11459 1919 11462
rect 3504 11456 3824 11457
rect 3504 11392 3512 11456
rect 3576 11392 3592 11456
rect 3656 11392 3672 11456
rect 3736 11392 3752 11456
rect 3816 11392 3824 11456
rect 3504 11391 3824 11392
rect 8626 11456 8946 11457
rect 8626 11392 8634 11456
rect 8698 11392 8714 11456
rect 8778 11392 8794 11456
rect 8858 11392 8874 11456
rect 8938 11392 8946 11456
rect 8626 11391 8946 11392
rect 13747 11456 14067 11457
rect 13747 11392 13755 11456
rect 13819 11392 13835 11456
rect 13899 11392 13915 11456
rect 13979 11392 13995 11456
rect 14059 11392 14067 11456
rect 13747 11391 14067 11392
rect 12525 11250 12591 11253
rect 16784 11250 17584 11280
rect 12525 11248 17584 11250
rect 12525 11192 12530 11248
rect 12586 11192 17584 11248
rect 12525 11190 17584 11192
rect 12525 11187 12591 11190
rect 16784 11160 17584 11190
rect 6065 10912 6385 10913
rect 6065 10848 6073 10912
rect 6137 10848 6153 10912
rect 6217 10848 6233 10912
rect 6297 10848 6313 10912
rect 6377 10848 6385 10912
rect 6065 10847 6385 10848
rect 11186 10912 11506 10913
rect 11186 10848 11194 10912
rect 11258 10848 11274 10912
rect 11338 10848 11354 10912
rect 11418 10848 11434 10912
rect 11498 10848 11506 10912
rect 11186 10847 11506 10848
rect 3504 10368 3824 10369
rect 3504 10304 3512 10368
rect 3576 10304 3592 10368
rect 3656 10304 3672 10368
rect 3736 10304 3752 10368
rect 3816 10304 3824 10368
rect 3504 10303 3824 10304
rect 8626 10368 8946 10369
rect 8626 10304 8634 10368
rect 8698 10304 8714 10368
rect 8778 10304 8794 10368
rect 8858 10304 8874 10368
rect 8938 10304 8946 10368
rect 8626 10303 8946 10304
rect 13747 10368 14067 10369
rect 13747 10304 13755 10368
rect 13819 10304 13835 10368
rect 13899 10304 13915 10368
rect 13979 10304 13995 10368
rect 14059 10304 14067 10368
rect 13747 10303 14067 10304
rect 6065 9824 6385 9825
rect 6065 9760 6073 9824
rect 6137 9760 6153 9824
rect 6217 9760 6233 9824
rect 6297 9760 6313 9824
rect 6377 9760 6385 9824
rect 6065 9759 6385 9760
rect 11186 9824 11506 9825
rect 11186 9760 11194 9824
rect 11258 9760 11274 9824
rect 11338 9760 11354 9824
rect 11418 9760 11434 9824
rect 11498 9760 11506 9824
rect 11186 9759 11506 9760
rect 3504 9280 3824 9281
rect 3504 9216 3512 9280
rect 3576 9216 3592 9280
rect 3656 9216 3672 9280
rect 3736 9216 3752 9280
rect 3816 9216 3824 9280
rect 3504 9215 3824 9216
rect 8626 9280 8946 9281
rect 8626 9216 8634 9280
rect 8698 9216 8714 9280
rect 8778 9216 8794 9280
rect 8858 9216 8874 9280
rect 8938 9216 8946 9280
rect 8626 9215 8946 9216
rect 13747 9280 14067 9281
rect 13747 9216 13755 9280
rect 13819 9216 13835 9280
rect 13899 9216 13915 9280
rect 13979 9216 13995 9280
rect 14059 9216 14067 9280
rect 13747 9215 14067 9216
rect 6065 8736 6385 8737
rect 6065 8672 6073 8736
rect 6137 8672 6153 8736
rect 6217 8672 6233 8736
rect 6297 8672 6313 8736
rect 6377 8672 6385 8736
rect 6065 8671 6385 8672
rect 11186 8736 11506 8737
rect 11186 8672 11194 8736
rect 11258 8672 11274 8736
rect 11338 8672 11354 8736
rect 11418 8672 11434 8736
rect 11498 8672 11506 8736
rect 11186 8671 11506 8672
rect 0 8530 800 8560
rect 2865 8530 2931 8533
rect 0 8528 2931 8530
rect 0 8472 2870 8528
rect 2926 8472 2931 8528
rect 0 8470 2931 8472
rect 0 8440 800 8470
rect 2865 8467 2931 8470
rect 15653 8258 15719 8261
rect 16784 8258 17584 8288
rect 15653 8256 17584 8258
rect 15653 8200 15658 8256
rect 15714 8200 17584 8256
rect 15653 8198 17584 8200
rect 15653 8195 15719 8198
rect 3504 8192 3824 8193
rect 3504 8128 3512 8192
rect 3576 8128 3592 8192
rect 3656 8128 3672 8192
rect 3736 8128 3752 8192
rect 3816 8128 3824 8192
rect 3504 8127 3824 8128
rect 8626 8192 8946 8193
rect 8626 8128 8634 8192
rect 8698 8128 8714 8192
rect 8778 8128 8794 8192
rect 8858 8128 8874 8192
rect 8938 8128 8946 8192
rect 8626 8127 8946 8128
rect 13747 8192 14067 8193
rect 13747 8128 13755 8192
rect 13819 8128 13835 8192
rect 13899 8128 13915 8192
rect 13979 8128 13995 8192
rect 14059 8128 14067 8192
rect 16784 8168 17584 8198
rect 13747 8127 14067 8128
rect 5349 7986 5415 7989
rect 12985 7986 13051 7989
rect 5349 7984 13051 7986
rect 5349 7928 5354 7984
rect 5410 7928 12990 7984
rect 13046 7928 13051 7984
rect 5349 7926 13051 7928
rect 5349 7923 5415 7926
rect 12985 7923 13051 7926
rect 6545 7850 6611 7853
rect 9857 7850 9923 7853
rect 6545 7848 9923 7850
rect 6545 7792 6550 7848
rect 6606 7792 9862 7848
rect 9918 7792 9923 7848
rect 6545 7790 9923 7792
rect 6545 7787 6611 7790
rect 9857 7787 9923 7790
rect 6637 7714 6703 7717
rect 8385 7714 8451 7717
rect 6637 7712 8451 7714
rect 6637 7656 6642 7712
rect 6698 7656 8390 7712
rect 8446 7656 8451 7712
rect 6637 7654 8451 7656
rect 6637 7651 6703 7654
rect 8385 7651 8451 7654
rect 6065 7648 6385 7649
rect 6065 7584 6073 7648
rect 6137 7584 6153 7648
rect 6217 7584 6233 7648
rect 6297 7584 6313 7648
rect 6377 7584 6385 7648
rect 6065 7583 6385 7584
rect 11186 7648 11506 7649
rect 11186 7584 11194 7648
rect 11258 7584 11274 7648
rect 11338 7584 11354 7648
rect 11418 7584 11434 7648
rect 11498 7584 11506 7648
rect 11186 7583 11506 7584
rect 7465 7578 7531 7581
rect 8293 7578 8359 7581
rect 7465 7576 8359 7578
rect 7465 7520 7470 7576
rect 7526 7520 8298 7576
rect 8354 7520 8359 7576
rect 7465 7518 8359 7520
rect 7465 7515 7531 7518
rect 8293 7515 8359 7518
rect 4613 7442 4679 7445
rect 11145 7442 11211 7445
rect 4613 7440 11211 7442
rect 4613 7384 4618 7440
rect 4674 7384 11150 7440
rect 11206 7384 11211 7440
rect 4613 7382 11211 7384
rect 4613 7379 4679 7382
rect 11145 7379 11211 7382
rect 4797 7306 4863 7309
rect 11513 7306 11579 7309
rect 4797 7304 11579 7306
rect 4797 7248 4802 7304
rect 4858 7248 11518 7304
rect 11574 7248 11579 7304
rect 4797 7246 11579 7248
rect 4797 7243 4863 7246
rect 11513 7243 11579 7246
rect 8017 7170 8083 7173
rect 8477 7170 8543 7173
rect 8017 7168 8543 7170
rect 8017 7112 8022 7168
rect 8078 7112 8482 7168
rect 8538 7112 8543 7168
rect 8017 7110 8543 7112
rect 8017 7107 8083 7110
rect 8477 7107 8543 7110
rect 3504 7104 3824 7105
rect 3504 7040 3512 7104
rect 3576 7040 3592 7104
rect 3656 7040 3672 7104
rect 3736 7040 3752 7104
rect 3816 7040 3824 7104
rect 3504 7039 3824 7040
rect 8626 7104 8946 7105
rect 8626 7040 8634 7104
rect 8698 7040 8714 7104
rect 8778 7040 8794 7104
rect 8858 7040 8874 7104
rect 8938 7040 8946 7104
rect 8626 7039 8946 7040
rect 13747 7104 14067 7105
rect 13747 7040 13755 7104
rect 13819 7040 13835 7104
rect 13899 7040 13915 7104
rect 13979 7040 13995 7104
rect 14059 7040 14067 7104
rect 13747 7039 14067 7040
rect 7005 7034 7071 7037
rect 8477 7034 8543 7037
rect 7005 7032 8543 7034
rect 7005 6976 7010 7032
rect 7066 6976 8482 7032
rect 8538 6976 8543 7032
rect 7005 6974 8543 6976
rect 7005 6971 7071 6974
rect 8477 6971 8543 6974
rect 10961 7034 11027 7037
rect 12709 7034 12775 7037
rect 10961 7032 12775 7034
rect 10961 6976 10966 7032
rect 11022 6976 12714 7032
rect 12770 6976 12775 7032
rect 10961 6974 12775 6976
rect 10961 6971 11027 6974
rect 12709 6971 12775 6974
rect 5349 6898 5415 6901
rect 9121 6898 9187 6901
rect 5349 6896 9187 6898
rect 5349 6840 5354 6896
rect 5410 6840 9126 6896
rect 9182 6840 9187 6896
rect 5349 6838 9187 6840
rect 5349 6835 5415 6838
rect 9121 6835 9187 6838
rect 11421 6898 11487 6901
rect 12893 6898 12959 6901
rect 11421 6896 12959 6898
rect 11421 6840 11426 6896
rect 11482 6840 12898 6896
rect 12954 6840 12959 6896
rect 11421 6838 12959 6840
rect 11421 6835 11487 6838
rect 12893 6835 12959 6838
rect 7465 6762 7531 6765
rect 7925 6762 7991 6765
rect 7465 6760 7991 6762
rect 7465 6704 7470 6760
rect 7526 6704 7930 6760
rect 7986 6704 7991 6760
rect 7465 6702 7991 6704
rect 7465 6699 7531 6702
rect 7925 6699 7991 6702
rect 9673 6762 9739 6765
rect 11789 6762 11855 6765
rect 9673 6760 11855 6762
rect 9673 6704 9678 6760
rect 9734 6704 11794 6760
rect 11850 6704 11855 6760
rect 9673 6702 11855 6704
rect 9673 6699 9739 6702
rect 11789 6699 11855 6702
rect 6637 6626 6703 6629
rect 7649 6626 7715 6629
rect 6637 6624 7715 6626
rect 6637 6568 6642 6624
rect 6698 6568 7654 6624
rect 7710 6568 7715 6624
rect 6637 6566 7715 6568
rect 6637 6563 6703 6566
rect 7649 6563 7715 6566
rect 6065 6560 6385 6561
rect 6065 6496 6073 6560
rect 6137 6496 6153 6560
rect 6217 6496 6233 6560
rect 6297 6496 6313 6560
rect 6377 6496 6385 6560
rect 6065 6495 6385 6496
rect 11186 6560 11506 6561
rect 11186 6496 11194 6560
rect 11258 6496 11274 6560
rect 11338 6496 11354 6560
rect 11418 6496 11434 6560
rect 11498 6496 11506 6560
rect 11186 6495 11506 6496
rect 7833 6490 7899 6493
rect 8150 6490 8156 6492
rect 7833 6488 8156 6490
rect 7833 6432 7838 6488
rect 7894 6432 8156 6488
rect 7833 6430 8156 6432
rect 7833 6427 7899 6430
rect 8150 6428 8156 6430
rect 8220 6428 8226 6492
rect 9765 6490 9831 6493
rect 10133 6490 10199 6493
rect 10317 6490 10383 6493
rect 9765 6488 10383 6490
rect 9765 6432 9770 6488
rect 9826 6432 10138 6488
rect 10194 6432 10322 6488
rect 10378 6432 10383 6488
rect 9765 6430 10383 6432
rect 9765 6427 9831 6430
rect 10133 6427 10199 6430
rect 10317 6427 10383 6430
rect 6453 6354 6519 6357
rect 10317 6354 10383 6357
rect 11789 6354 11855 6357
rect 6453 6352 11855 6354
rect 6453 6296 6458 6352
rect 6514 6296 10322 6352
rect 10378 6296 11794 6352
rect 11850 6296 11855 6352
rect 6453 6294 11855 6296
rect 6453 6291 6519 6294
rect 10317 6291 10383 6294
rect 11789 6291 11855 6294
rect 9765 6218 9831 6221
rect 13721 6218 13787 6221
rect 9765 6216 13787 6218
rect 9765 6160 9770 6216
rect 9826 6160 13726 6216
rect 13782 6160 13787 6216
rect 9765 6158 13787 6160
rect 9765 6155 9831 6158
rect 13721 6155 13787 6158
rect 3504 6016 3824 6017
rect 3504 5952 3512 6016
rect 3576 5952 3592 6016
rect 3656 5952 3672 6016
rect 3736 5952 3752 6016
rect 3816 5952 3824 6016
rect 3504 5951 3824 5952
rect 8626 6016 8946 6017
rect 8626 5952 8634 6016
rect 8698 5952 8714 6016
rect 8778 5952 8794 6016
rect 8858 5952 8874 6016
rect 8938 5952 8946 6016
rect 8626 5951 8946 5952
rect 13747 6016 14067 6017
rect 13747 5952 13755 6016
rect 13819 5952 13835 6016
rect 13899 5952 13915 6016
rect 13979 5952 13995 6016
rect 14059 5952 14067 6016
rect 13747 5951 14067 5952
rect 5901 5946 5967 5949
rect 8201 5946 8267 5949
rect 5901 5944 8267 5946
rect 5901 5888 5906 5944
rect 5962 5888 8206 5944
rect 8262 5888 8267 5944
rect 5901 5886 8267 5888
rect 5901 5883 5967 5886
rect 8201 5883 8267 5886
rect 0 5810 800 5840
rect 1393 5810 1459 5813
rect 0 5808 1459 5810
rect 0 5752 1398 5808
rect 1454 5752 1459 5808
rect 0 5750 1459 5752
rect 0 5720 800 5750
rect 1393 5747 1459 5750
rect 2497 5810 2563 5813
rect 2773 5810 2839 5813
rect 2497 5808 2839 5810
rect 2497 5752 2502 5808
rect 2558 5752 2778 5808
rect 2834 5752 2839 5808
rect 2497 5750 2839 5752
rect 2497 5747 2563 5750
rect 2773 5747 2839 5750
rect 14273 5538 14339 5541
rect 16784 5538 17584 5568
rect 14273 5536 17584 5538
rect 14273 5480 14278 5536
rect 14334 5480 17584 5536
rect 14273 5478 17584 5480
rect 14273 5475 14339 5478
rect 6065 5472 6385 5473
rect 6065 5408 6073 5472
rect 6137 5408 6153 5472
rect 6217 5408 6233 5472
rect 6297 5408 6313 5472
rect 6377 5408 6385 5472
rect 6065 5407 6385 5408
rect 11186 5472 11506 5473
rect 11186 5408 11194 5472
rect 11258 5408 11274 5472
rect 11338 5408 11354 5472
rect 11418 5408 11434 5472
rect 11498 5408 11506 5472
rect 16784 5448 17584 5478
rect 11186 5407 11506 5408
rect 3504 4928 3824 4929
rect 3504 4864 3512 4928
rect 3576 4864 3592 4928
rect 3656 4864 3672 4928
rect 3736 4864 3752 4928
rect 3816 4864 3824 4928
rect 3504 4863 3824 4864
rect 8626 4928 8946 4929
rect 8626 4864 8634 4928
rect 8698 4864 8714 4928
rect 8778 4864 8794 4928
rect 8858 4864 8874 4928
rect 8938 4864 8946 4928
rect 8626 4863 8946 4864
rect 13747 4928 14067 4929
rect 13747 4864 13755 4928
rect 13819 4864 13835 4928
rect 13899 4864 13915 4928
rect 13979 4864 13995 4928
rect 14059 4864 14067 4928
rect 13747 4863 14067 4864
rect 6065 4384 6385 4385
rect 6065 4320 6073 4384
rect 6137 4320 6153 4384
rect 6217 4320 6233 4384
rect 6297 4320 6313 4384
rect 6377 4320 6385 4384
rect 6065 4319 6385 4320
rect 11186 4384 11506 4385
rect 11186 4320 11194 4384
rect 11258 4320 11274 4384
rect 11338 4320 11354 4384
rect 11418 4320 11434 4384
rect 11498 4320 11506 4384
rect 11186 4319 11506 4320
rect 7281 4314 7347 4317
rect 8385 4314 8451 4317
rect 9213 4314 9279 4317
rect 7281 4312 9279 4314
rect 7281 4256 7286 4312
rect 7342 4256 8390 4312
rect 8446 4256 9218 4312
rect 9274 4256 9279 4312
rect 7281 4254 9279 4256
rect 7281 4251 7347 4254
rect 8385 4251 8451 4254
rect 9213 4251 9279 4254
rect 8201 4178 8267 4181
rect 9397 4178 9463 4181
rect 8201 4176 9463 4178
rect 8201 4120 8206 4176
rect 8262 4120 9402 4176
rect 9458 4120 9463 4176
rect 8201 4118 9463 4120
rect 8201 4115 8267 4118
rect 9397 4115 9463 4118
rect 7097 4042 7163 4045
rect 8293 4042 8359 4045
rect 7097 4040 8359 4042
rect 7097 3984 7102 4040
rect 7158 3984 8298 4040
rect 8354 3984 8359 4040
rect 7097 3982 8359 3984
rect 7097 3979 7163 3982
rect 8293 3979 8359 3982
rect 3504 3840 3824 3841
rect 3504 3776 3512 3840
rect 3576 3776 3592 3840
rect 3656 3776 3672 3840
rect 3736 3776 3752 3840
rect 3816 3776 3824 3840
rect 3504 3775 3824 3776
rect 8626 3840 8946 3841
rect 8626 3776 8634 3840
rect 8698 3776 8714 3840
rect 8778 3776 8794 3840
rect 8858 3776 8874 3840
rect 8938 3776 8946 3840
rect 8626 3775 8946 3776
rect 13747 3840 14067 3841
rect 13747 3776 13755 3840
rect 13819 3776 13835 3840
rect 13899 3776 13915 3840
rect 13979 3776 13995 3840
rect 14059 3776 14067 3840
rect 13747 3775 14067 3776
rect 3877 3634 3943 3637
rect 7741 3634 7807 3637
rect 3877 3632 7807 3634
rect 3877 3576 3882 3632
rect 3938 3576 7746 3632
rect 7802 3576 7807 3632
rect 3877 3574 7807 3576
rect 3877 3571 3943 3574
rect 7741 3571 7807 3574
rect 2681 3498 2747 3501
rect 6085 3498 6151 3501
rect 2681 3496 6151 3498
rect 2681 3440 2686 3496
rect 2742 3440 6090 3496
rect 6146 3440 6151 3496
rect 2681 3438 6151 3440
rect 2681 3435 2747 3438
rect 6085 3435 6151 3438
rect 7189 3498 7255 3501
rect 8293 3498 8359 3501
rect 7189 3496 8359 3498
rect 7189 3440 7194 3496
rect 7250 3440 8298 3496
rect 8354 3440 8359 3496
rect 7189 3438 8359 3440
rect 7189 3435 7255 3438
rect 8293 3435 8359 3438
rect 6065 3296 6385 3297
rect 6065 3232 6073 3296
rect 6137 3232 6153 3296
rect 6217 3232 6233 3296
rect 6297 3232 6313 3296
rect 6377 3232 6385 3296
rect 6065 3231 6385 3232
rect 11186 3296 11506 3297
rect 11186 3232 11194 3296
rect 11258 3232 11274 3296
rect 11338 3232 11354 3296
rect 11418 3232 11434 3296
rect 11498 3232 11506 3296
rect 11186 3231 11506 3232
rect 2589 3226 2655 3229
rect 5625 3226 5691 3229
rect 2589 3224 5691 3226
rect 2589 3168 2594 3224
rect 2650 3168 5630 3224
rect 5686 3168 5691 3224
rect 2589 3166 5691 3168
rect 2589 3163 2655 3166
rect 5625 3163 5691 3166
rect 1577 3090 1643 3093
rect 7097 3090 7163 3093
rect 1577 3088 7163 3090
rect 1577 3032 1582 3088
rect 1638 3032 7102 3088
rect 7158 3032 7163 3088
rect 1577 3030 7163 3032
rect 1577 3027 1643 3030
rect 7097 3027 7163 3030
rect 7281 3090 7347 3093
rect 8753 3090 8819 3093
rect 7281 3088 8819 3090
rect 7281 3032 7286 3088
rect 7342 3032 8758 3088
rect 8814 3032 8819 3088
rect 7281 3030 8819 3032
rect 7281 3027 7347 3030
rect 8753 3027 8819 3030
rect 4429 2954 4495 2957
rect 7005 2954 7071 2957
rect 4429 2952 7071 2954
rect 4429 2896 4434 2952
rect 4490 2896 7010 2952
rect 7066 2896 7071 2952
rect 4429 2894 7071 2896
rect 4429 2891 4495 2894
rect 7005 2891 7071 2894
rect 8150 2892 8156 2956
rect 8220 2954 8226 2956
rect 10041 2954 10107 2957
rect 8220 2952 10107 2954
rect 8220 2896 10046 2952
rect 10102 2896 10107 2952
rect 8220 2894 10107 2896
rect 8220 2892 8226 2894
rect 10041 2891 10107 2894
rect 0 2818 800 2848
rect 2773 2818 2839 2821
rect 0 2816 2839 2818
rect 0 2760 2778 2816
rect 2834 2760 2839 2816
rect 0 2758 2839 2760
rect 0 2728 800 2758
rect 2773 2755 2839 2758
rect 3504 2752 3824 2753
rect 3504 2688 3512 2752
rect 3576 2688 3592 2752
rect 3656 2688 3672 2752
rect 3736 2688 3752 2752
rect 3816 2688 3824 2752
rect 3504 2687 3824 2688
rect 8626 2752 8946 2753
rect 8626 2688 8634 2752
rect 8698 2688 8714 2752
rect 8778 2688 8794 2752
rect 8858 2688 8874 2752
rect 8938 2688 8946 2752
rect 8626 2687 8946 2688
rect 13747 2752 14067 2753
rect 13747 2688 13755 2752
rect 13819 2688 13835 2752
rect 13899 2688 13915 2752
rect 13979 2688 13995 2752
rect 14059 2688 14067 2752
rect 13747 2687 14067 2688
rect 15745 2546 15811 2549
rect 16784 2546 17584 2576
rect 15745 2544 17584 2546
rect 15745 2488 15750 2544
rect 15806 2488 17584 2544
rect 15745 2486 17584 2488
rect 15745 2483 15811 2486
rect 16784 2456 17584 2486
rect 6065 2208 6385 2209
rect 6065 2144 6073 2208
rect 6137 2144 6153 2208
rect 6217 2144 6233 2208
rect 6297 2144 6313 2208
rect 6377 2144 6385 2208
rect 6065 2143 6385 2144
rect 11186 2208 11506 2209
rect 11186 2144 11194 2208
rect 11258 2144 11274 2208
rect 11338 2144 11354 2208
rect 11418 2144 11434 2208
rect 11498 2144 11506 2208
rect 11186 2143 11506 2144
<< via3 >>
rect 6073 17436 6137 17440
rect 6073 17380 6077 17436
rect 6077 17380 6133 17436
rect 6133 17380 6137 17436
rect 6073 17376 6137 17380
rect 6153 17436 6217 17440
rect 6153 17380 6157 17436
rect 6157 17380 6213 17436
rect 6213 17380 6217 17436
rect 6153 17376 6217 17380
rect 6233 17436 6297 17440
rect 6233 17380 6237 17436
rect 6237 17380 6293 17436
rect 6293 17380 6297 17436
rect 6233 17376 6297 17380
rect 6313 17436 6377 17440
rect 6313 17380 6317 17436
rect 6317 17380 6373 17436
rect 6373 17380 6377 17436
rect 6313 17376 6377 17380
rect 11194 17436 11258 17440
rect 11194 17380 11198 17436
rect 11198 17380 11254 17436
rect 11254 17380 11258 17436
rect 11194 17376 11258 17380
rect 11274 17436 11338 17440
rect 11274 17380 11278 17436
rect 11278 17380 11334 17436
rect 11334 17380 11338 17436
rect 11274 17376 11338 17380
rect 11354 17436 11418 17440
rect 11354 17380 11358 17436
rect 11358 17380 11414 17436
rect 11414 17380 11418 17436
rect 11354 17376 11418 17380
rect 11434 17436 11498 17440
rect 11434 17380 11438 17436
rect 11438 17380 11494 17436
rect 11494 17380 11498 17436
rect 11434 17376 11498 17380
rect 3512 16892 3576 16896
rect 3512 16836 3516 16892
rect 3516 16836 3572 16892
rect 3572 16836 3576 16892
rect 3512 16832 3576 16836
rect 3592 16892 3656 16896
rect 3592 16836 3596 16892
rect 3596 16836 3652 16892
rect 3652 16836 3656 16892
rect 3592 16832 3656 16836
rect 3672 16892 3736 16896
rect 3672 16836 3676 16892
rect 3676 16836 3732 16892
rect 3732 16836 3736 16892
rect 3672 16832 3736 16836
rect 3752 16892 3816 16896
rect 3752 16836 3756 16892
rect 3756 16836 3812 16892
rect 3812 16836 3816 16892
rect 3752 16832 3816 16836
rect 8634 16892 8698 16896
rect 8634 16836 8638 16892
rect 8638 16836 8694 16892
rect 8694 16836 8698 16892
rect 8634 16832 8698 16836
rect 8714 16892 8778 16896
rect 8714 16836 8718 16892
rect 8718 16836 8774 16892
rect 8774 16836 8778 16892
rect 8714 16832 8778 16836
rect 8794 16892 8858 16896
rect 8794 16836 8798 16892
rect 8798 16836 8854 16892
rect 8854 16836 8858 16892
rect 8794 16832 8858 16836
rect 8874 16892 8938 16896
rect 8874 16836 8878 16892
rect 8878 16836 8934 16892
rect 8934 16836 8938 16892
rect 8874 16832 8938 16836
rect 13755 16892 13819 16896
rect 13755 16836 13759 16892
rect 13759 16836 13815 16892
rect 13815 16836 13819 16892
rect 13755 16832 13819 16836
rect 13835 16892 13899 16896
rect 13835 16836 13839 16892
rect 13839 16836 13895 16892
rect 13895 16836 13899 16892
rect 13835 16832 13899 16836
rect 13915 16892 13979 16896
rect 13915 16836 13919 16892
rect 13919 16836 13975 16892
rect 13975 16836 13979 16892
rect 13915 16832 13979 16836
rect 13995 16892 14059 16896
rect 13995 16836 13999 16892
rect 13999 16836 14055 16892
rect 14055 16836 14059 16892
rect 13995 16832 14059 16836
rect 6073 16348 6137 16352
rect 6073 16292 6077 16348
rect 6077 16292 6133 16348
rect 6133 16292 6137 16348
rect 6073 16288 6137 16292
rect 6153 16348 6217 16352
rect 6153 16292 6157 16348
rect 6157 16292 6213 16348
rect 6213 16292 6217 16348
rect 6153 16288 6217 16292
rect 6233 16348 6297 16352
rect 6233 16292 6237 16348
rect 6237 16292 6293 16348
rect 6293 16292 6297 16348
rect 6233 16288 6297 16292
rect 6313 16348 6377 16352
rect 6313 16292 6317 16348
rect 6317 16292 6373 16348
rect 6373 16292 6377 16348
rect 6313 16288 6377 16292
rect 11194 16348 11258 16352
rect 11194 16292 11198 16348
rect 11198 16292 11254 16348
rect 11254 16292 11258 16348
rect 11194 16288 11258 16292
rect 11274 16348 11338 16352
rect 11274 16292 11278 16348
rect 11278 16292 11334 16348
rect 11334 16292 11338 16348
rect 11274 16288 11338 16292
rect 11354 16348 11418 16352
rect 11354 16292 11358 16348
rect 11358 16292 11414 16348
rect 11414 16292 11418 16348
rect 11354 16288 11418 16292
rect 11434 16348 11498 16352
rect 11434 16292 11438 16348
rect 11438 16292 11494 16348
rect 11494 16292 11498 16348
rect 11434 16288 11498 16292
rect 3512 15804 3576 15808
rect 3512 15748 3516 15804
rect 3516 15748 3572 15804
rect 3572 15748 3576 15804
rect 3512 15744 3576 15748
rect 3592 15804 3656 15808
rect 3592 15748 3596 15804
rect 3596 15748 3652 15804
rect 3652 15748 3656 15804
rect 3592 15744 3656 15748
rect 3672 15804 3736 15808
rect 3672 15748 3676 15804
rect 3676 15748 3732 15804
rect 3732 15748 3736 15804
rect 3672 15744 3736 15748
rect 3752 15804 3816 15808
rect 3752 15748 3756 15804
rect 3756 15748 3812 15804
rect 3812 15748 3816 15804
rect 3752 15744 3816 15748
rect 8634 15804 8698 15808
rect 8634 15748 8638 15804
rect 8638 15748 8694 15804
rect 8694 15748 8698 15804
rect 8634 15744 8698 15748
rect 8714 15804 8778 15808
rect 8714 15748 8718 15804
rect 8718 15748 8774 15804
rect 8774 15748 8778 15804
rect 8714 15744 8778 15748
rect 8794 15804 8858 15808
rect 8794 15748 8798 15804
rect 8798 15748 8854 15804
rect 8854 15748 8858 15804
rect 8794 15744 8858 15748
rect 8874 15804 8938 15808
rect 8874 15748 8878 15804
rect 8878 15748 8934 15804
rect 8934 15748 8938 15804
rect 8874 15744 8938 15748
rect 13755 15804 13819 15808
rect 13755 15748 13759 15804
rect 13759 15748 13815 15804
rect 13815 15748 13819 15804
rect 13755 15744 13819 15748
rect 13835 15804 13899 15808
rect 13835 15748 13839 15804
rect 13839 15748 13895 15804
rect 13895 15748 13899 15804
rect 13835 15744 13899 15748
rect 13915 15804 13979 15808
rect 13915 15748 13919 15804
rect 13919 15748 13975 15804
rect 13975 15748 13979 15804
rect 13915 15744 13979 15748
rect 13995 15804 14059 15808
rect 13995 15748 13999 15804
rect 13999 15748 14055 15804
rect 14055 15748 14059 15804
rect 13995 15744 14059 15748
rect 6073 15260 6137 15264
rect 6073 15204 6077 15260
rect 6077 15204 6133 15260
rect 6133 15204 6137 15260
rect 6073 15200 6137 15204
rect 6153 15260 6217 15264
rect 6153 15204 6157 15260
rect 6157 15204 6213 15260
rect 6213 15204 6217 15260
rect 6153 15200 6217 15204
rect 6233 15260 6297 15264
rect 6233 15204 6237 15260
rect 6237 15204 6293 15260
rect 6293 15204 6297 15260
rect 6233 15200 6297 15204
rect 6313 15260 6377 15264
rect 6313 15204 6317 15260
rect 6317 15204 6373 15260
rect 6373 15204 6377 15260
rect 6313 15200 6377 15204
rect 11194 15260 11258 15264
rect 11194 15204 11198 15260
rect 11198 15204 11254 15260
rect 11254 15204 11258 15260
rect 11194 15200 11258 15204
rect 11274 15260 11338 15264
rect 11274 15204 11278 15260
rect 11278 15204 11334 15260
rect 11334 15204 11338 15260
rect 11274 15200 11338 15204
rect 11354 15260 11418 15264
rect 11354 15204 11358 15260
rect 11358 15204 11414 15260
rect 11414 15204 11418 15260
rect 11354 15200 11418 15204
rect 11434 15260 11498 15264
rect 11434 15204 11438 15260
rect 11438 15204 11494 15260
rect 11494 15204 11498 15260
rect 11434 15200 11498 15204
rect 3512 14716 3576 14720
rect 3512 14660 3516 14716
rect 3516 14660 3572 14716
rect 3572 14660 3576 14716
rect 3512 14656 3576 14660
rect 3592 14716 3656 14720
rect 3592 14660 3596 14716
rect 3596 14660 3652 14716
rect 3652 14660 3656 14716
rect 3592 14656 3656 14660
rect 3672 14716 3736 14720
rect 3672 14660 3676 14716
rect 3676 14660 3732 14716
rect 3732 14660 3736 14716
rect 3672 14656 3736 14660
rect 3752 14716 3816 14720
rect 3752 14660 3756 14716
rect 3756 14660 3812 14716
rect 3812 14660 3816 14716
rect 3752 14656 3816 14660
rect 8634 14716 8698 14720
rect 8634 14660 8638 14716
rect 8638 14660 8694 14716
rect 8694 14660 8698 14716
rect 8634 14656 8698 14660
rect 8714 14716 8778 14720
rect 8714 14660 8718 14716
rect 8718 14660 8774 14716
rect 8774 14660 8778 14716
rect 8714 14656 8778 14660
rect 8794 14716 8858 14720
rect 8794 14660 8798 14716
rect 8798 14660 8854 14716
rect 8854 14660 8858 14716
rect 8794 14656 8858 14660
rect 8874 14716 8938 14720
rect 8874 14660 8878 14716
rect 8878 14660 8934 14716
rect 8934 14660 8938 14716
rect 8874 14656 8938 14660
rect 13755 14716 13819 14720
rect 13755 14660 13759 14716
rect 13759 14660 13815 14716
rect 13815 14660 13819 14716
rect 13755 14656 13819 14660
rect 13835 14716 13899 14720
rect 13835 14660 13839 14716
rect 13839 14660 13895 14716
rect 13895 14660 13899 14716
rect 13835 14656 13899 14660
rect 13915 14716 13979 14720
rect 13915 14660 13919 14716
rect 13919 14660 13975 14716
rect 13975 14660 13979 14716
rect 13915 14656 13979 14660
rect 13995 14716 14059 14720
rect 13995 14660 13999 14716
rect 13999 14660 14055 14716
rect 14055 14660 14059 14716
rect 13995 14656 14059 14660
rect 6073 14172 6137 14176
rect 6073 14116 6077 14172
rect 6077 14116 6133 14172
rect 6133 14116 6137 14172
rect 6073 14112 6137 14116
rect 6153 14172 6217 14176
rect 6153 14116 6157 14172
rect 6157 14116 6213 14172
rect 6213 14116 6217 14172
rect 6153 14112 6217 14116
rect 6233 14172 6297 14176
rect 6233 14116 6237 14172
rect 6237 14116 6293 14172
rect 6293 14116 6297 14172
rect 6233 14112 6297 14116
rect 6313 14172 6377 14176
rect 6313 14116 6317 14172
rect 6317 14116 6373 14172
rect 6373 14116 6377 14172
rect 6313 14112 6377 14116
rect 11194 14172 11258 14176
rect 11194 14116 11198 14172
rect 11198 14116 11254 14172
rect 11254 14116 11258 14172
rect 11194 14112 11258 14116
rect 11274 14172 11338 14176
rect 11274 14116 11278 14172
rect 11278 14116 11334 14172
rect 11334 14116 11338 14172
rect 11274 14112 11338 14116
rect 11354 14172 11418 14176
rect 11354 14116 11358 14172
rect 11358 14116 11414 14172
rect 11414 14116 11418 14172
rect 11354 14112 11418 14116
rect 11434 14172 11498 14176
rect 11434 14116 11438 14172
rect 11438 14116 11494 14172
rect 11494 14116 11498 14172
rect 11434 14112 11498 14116
rect 3512 13628 3576 13632
rect 3512 13572 3516 13628
rect 3516 13572 3572 13628
rect 3572 13572 3576 13628
rect 3512 13568 3576 13572
rect 3592 13628 3656 13632
rect 3592 13572 3596 13628
rect 3596 13572 3652 13628
rect 3652 13572 3656 13628
rect 3592 13568 3656 13572
rect 3672 13628 3736 13632
rect 3672 13572 3676 13628
rect 3676 13572 3732 13628
rect 3732 13572 3736 13628
rect 3672 13568 3736 13572
rect 3752 13628 3816 13632
rect 3752 13572 3756 13628
rect 3756 13572 3812 13628
rect 3812 13572 3816 13628
rect 3752 13568 3816 13572
rect 8634 13628 8698 13632
rect 8634 13572 8638 13628
rect 8638 13572 8694 13628
rect 8694 13572 8698 13628
rect 8634 13568 8698 13572
rect 8714 13628 8778 13632
rect 8714 13572 8718 13628
rect 8718 13572 8774 13628
rect 8774 13572 8778 13628
rect 8714 13568 8778 13572
rect 8794 13628 8858 13632
rect 8794 13572 8798 13628
rect 8798 13572 8854 13628
rect 8854 13572 8858 13628
rect 8794 13568 8858 13572
rect 8874 13628 8938 13632
rect 8874 13572 8878 13628
rect 8878 13572 8934 13628
rect 8934 13572 8938 13628
rect 8874 13568 8938 13572
rect 13755 13628 13819 13632
rect 13755 13572 13759 13628
rect 13759 13572 13815 13628
rect 13815 13572 13819 13628
rect 13755 13568 13819 13572
rect 13835 13628 13899 13632
rect 13835 13572 13839 13628
rect 13839 13572 13895 13628
rect 13895 13572 13899 13628
rect 13835 13568 13899 13572
rect 13915 13628 13979 13632
rect 13915 13572 13919 13628
rect 13919 13572 13975 13628
rect 13975 13572 13979 13628
rect 13915 13568 13979 13572
rect 13995 13628 14059 13632
rect 13995 13572 13999 13628
rect 13999 13572 14055 13628
rect 14055 13572 14059 13628
rect 13995 13568 14059 13572
rect 6073 13084 6137 13088
rect 6073 13028 6077 13084
rect 6077 13028 6133 13084
rect 6133 13028 6137 13084
rect 6073 13024 6137 13028
rect 6153 13084 6217 13088
rect 6153 13028 6157 13084
rect 6157 13028 6213 13084
rect 6213 13028 6217 13084
rect 6153 13024 6217 13028
rect 6233 13084 6297 13088
rect 6233 13028 6237 13084
rect 6237 13028 6293 13084
rect 6293 13028 6297 13084
rect 6233 13024 6297 13028
rect 6313 13084 6377 13088
rect 6313 13028 6317 13084
rect 6317 13028 6373 13084
rect 6373 13028 6377 13084
rect 6313 13024 6377 13028
rect 11194 13084 11258 13088
rect 11194 13028 11198 13084
rect 11198 13028 11254 13084
rect 11254 13028 11258 13084
rect 11194 13024 11258 13028
rect 11274 13084 11338 13088
rect 11274 13028 11278 13084
rect 11278 13028 11334 13084
rect 11334 13028 11338 13084
rect 11274 13024 11338 13028
rect 11354 13084 11418 13088
rect 11354 13028 11358 13084
rect 11358 13028 11414 13084
rect 11414 13028 11418 13084
rect 11354 13024 11418 13028
rect 11434 13084 11498 13088
rect 11434 13028 11438 13084
rect 11438 13028 11494 13084
rect 11494 13028 11498 13084
rect 11434 13024 11498 13028
rect 3512 12540 3576 12544
rect 3512 12484 3516 12540
rect 3516 12484 3572 12540
rect 3572 12484 3576 12540
rect 3512 12480 3576 12484
rect 3592 12540 3656 12544
rect 3592 12484 3596 12540
rect 3596 12484 3652 12540
rect 3652 12484 3656 12540
rect 3592 12480 3656 12484
rect 3672 12540 3736 12544
rect 3672 12484 3676 12540
rect 3676 12484 3732 12540
rect 3732 12484 3736 12540
rect 3672 12480 3736 12484
rect 3752 12540 3816 12544
rect 3752 12484 3756 12540
rect 3756 12484 3812 12540
rect 3812 12484 3816 12540
rect 3752 12480 3816 12484
rect 8634 12540 8698 12544
rect 8634 12484 8638 12540
rect 8638 12484 8694 12540
rect 8694 12484 8698 12540
rect 8634 12480 8698 12484
rect 8714 12540 8778 12544
rect 8714 12484 8718 12540
rect 8718 12484 8774 12540
rect 8774 12484 8778 12540
rect 8714 12480 8778 12484
rect 8794 12540 8858 12544
rect 8794 12484 8798 12540
rect 8798 12484 8854 12540
rect 8854 12484 8858 12540
rect 8794 12480 8858 12484
rect 8874 12540 8938 12544
rect 8874 12484 8878 12540
rect 8878 12484 8934 12540
rect 8934 12484 8938 12540
rect 8874 12480 8938 12484
rect 13755 12540 13819 12544
rect 13755 12484 13759 12540
rect 13759 12484 13815 12540
rect 13815 12484 13819 12540
rect 13755 12480 13819 12484
rect 13835 12540 13899 12544
rect 13835 12484 13839 12540
rect 13839 12484 13895 12540
rect 13895 12484 13899 12540
rect 13835 12480 13899 12484
rect 13915 12540 13979 12544
rect 13915 12484 13919 12540
rect 13919 12484 13975 12540
rect 13975 12484 13979 12540
rect 13915 12480 13979 12484
rect 13995 12540 14059 12544
rect 13995 12484 13999 12540
rect 13999 12484 14055 12540
rect 14055 12484 14059 12540
rect 13995 12480 14059 12484
rect 6073 11996 6137 12000
rect 6073 11940 6077 11996
rect 6077 11940 6133 11996
rect 6133 11940 6137 11996
rect 6073 11936 6137 11940
rect 6153 11996 6217 12000
rect 6153 11940 6157 11996
rect 6157 11940 6213 11996
rect 6213 11940 6217 11996
rect 6153 11936 6217 11940
rect 6233 11996 6297 12000
rect 6233 11940 6237 11996
rect 6237 11940 6293 11996
rect 6293 11940 6297 11996
rect 6233 11936 6297 11940
rect 6313 11996 6377 12000
rect 6313 11940 6317 11996
rect 6317 11940 6373 11996
rect 6373 11940 6377 11996
rect 6313 11936 6377 11940
rect 11194 11996 11258 12000
rect 11194 11940 11198 11996
rect 11198 11940 11254 11996
rect 11254 11940 11258 11996
rect 11194 11936 11258 11940
rect 11274 11996 11338 12000
rect 11274 11940 11278 11996
rect 11278 11940 11334 11996
rect 11334 11940 11338 11996
rect 11274 11936 11338 11940
rect 11354 11996 11418 12000
rect 11354 11940 11358 11996
rect 11358 11940 11414 11996
rect 11414 11940 11418 11996
rect 11354 11936 11418 11940
rect 11434 11996 11498 12000
rect 11434 11940 11438 11996
rect 11438 11940 11494 11996
rect 11494 11940 11498 11996
rect 11434 11936 11498 11940
rect 3512 11452 3576 11456
rect 3512 11396 3516 11452
rect 3516 11396 3572 11452
rect 3572 11396 3576 11452
rect 3512 11392 3576 11396
rect 3592 11452 3656 11456
rect 3592 11396 3596 11452
rect 3596 11396 3652 11452
rect 3652 11396 3656 11452
rect 3592 11392 3656 11396
rect 3672 11452 3736 11456
rect 3672 11396 3676 11452
rect 3676 11396 3732 11452
rect 3732 11396 3736 11452
rect 3672 11392 3736 11396
rect 3752 11452 3816 11456
rect 3752 11396 3756 11452
rect 3756 11396 3812 11452
rect 3812 11396 3816 11452
rect 3752 11392 3816 11396
rect 8634 11452 8698 11456
rect 8634 11396 8638 11452
rect 8638 11396 8694 11452
rect 8694 11396 8698 11452
rect 8634 11392 8698 11396
rect 8714 11452 8778 11456
rect 8714 11396 8718 11452
rect 8718 11396 8774 11452
rect 8774 11396 8778 11452
rect 8714 11392 8778 11396
rect 8794 11452 8858 11456
rect 8794 11396 8798 11452
rect 8798 11396 8854 11452
rect 8854 11396 8858 11452
rect 8794 11392 8858 11396
rect 8874 11452 8938 11456
rect 8874 11396 8878 11452
rect 8878 11396 8934 11452
rect 8934 11396 8938 11452
rect 8874 11392 8938 11396
rect 13755 11452 13819 11456
rect 13755 11396 13759 11452
rect 13759 11396 13815 11452
rect 13815 11396 13819 11452
rect 13755 11392 13819 11396
rect 13835 11452 13899 11456
rect 13835 11396 13839 11452
rect 13839 11396 13895 11452
rect 13895 11396 13899 11452
rect 13835 11392 13899 11396
rect 13915 11452 13979 11456
rect 13915 11396 13919 11452
rect 13919 11396 13975 11452
rect 13975 11396 13979 11452
rect 13915 11392 13979 11396
rect 13995 11452 14059 11456
rect 13995 11396 13999 11452
rect 13999 11396 14055 11452
rect 14055 11396 14059 11452
rect 13995 11392 14059 11396
rect 6073 10908 6137 10912
rect 6073 10852 6077 10908
rect 6077 10852 6133 10908
rect 6133 10852 6137 10908
rect 6073 10848 6137 10852
rect 6153 10908 6217 10912
rect 6153 10852 6157 10908
rect 6157 10852 6213 10908
rect 6213 10852 6217 10908
rect 6153 10848 6217 10852
rect 6233 10908 6297 10912
rect 6233 10852 6237 10908
rect 6237 10852 6293 10908
rect 6293 10852 6297 10908
rect 6233 10848 6297 10852
rect 6313 10908 6377 10912
rect 6313 10852 6317 10908
rect 6317 10852 6373 10908
rect 6373 10852 6377 10908
rect 6313 10848 6377 10852
rect 11194 10908 11258 10912
rect 11194 10852 11198 10908
rect 11198 10852 11254 10908
rect 11254 10852 11258 10908
rect 11194 10848 11258 10852
rect 11274 10908 11338 10912
rect 11274 10852 11278 10908
rect 11278 10852 11334 10908
rect 11334 10852 11338 10908
rect 11274 10848 11338 10852
rect 11354 10908 11418 10912
rect 11354 10852 11358 10908
rect 11358 10852 11414 10908
rect 11414 10852 11418 10908
rect 11354 10848 11418 10852
rect 11434 10908 11498 10912
rect 11434 10852 11438 10908
rect 11438 10852 11494 10908
rect 11494 10852 11498 10908
rect 11434 10848 11498 10852
rect 3512 10364 3576 10368
rect 3512 10308 3516 10364
rect 3516 10308 3572 10364
rect 3572 10308 3576 10364
rect 3512 10304 3576 10308
rect 3592 10364 3656 10368
rect 3592 10308 3596 10364
rect 3596 10308 3652 10364
rect 3652 10308 3656 10364
rect 3592 10304 3656 10308
rect 3672 10364 3736 10368
rect 3672 10308 3676 10364
rect 3676 10308 3732 10364
rect 3732 10308 3736 10364
rect 3672 10304 3736 10308
rect 3752 10364 3816 10368
rect 3752 10308 3756 10364
rect 3756 10308 3812 10364
rect 3812 10308 3816 10364
rect 3752 10304 3816 10308
rect 8634 10364 8698 10368
rect 8634 10308 8638 10364
rect 8638 10308 8694 10364
rect 8694 10308 8698 10364
rect 8634 10304 8698 10308
rect 8714 10364 8778 10368
rect 8714 10308 8718 10364
rect 8718 10308 8774 10364
rect 8774 10308 8778 10364
rect 8714 10304 8778 10308
rect 8794 10364 8858 10368
rect 8794 10308 8798 10364
rect 8798 10308 8854 10364
rect 8854 10308 8858 10364
rect 8794 10304 8858 10308
rect 8874 10364 8938 10368
rect 8874 10308 8878 10364
rect 8878 10308 8934 10364
rect 8934 10308 8938 10364
rect 8874 10304 8938 10308
rect 13755 10364 13819 10368
rect 13755 10308 13759 10364
rect 13759 10308 13815 10364
rect 13815 10308 13819 10364
rect 13755 10304 13819 10308
rect 13835 10364 13899 10368
rect 13835 10308 13839 10364
rect 13839 10308 13895 10364
rect 13895 10308 13899 10364
rect 13835 10304 13899 10308
rect 13915 10364 13979 10368
rect 13915 10308 13919 10364
rect 13919 10308 13975 10364
rect 13975 10308 13979 10364
rect 13915 10304 13979 10308
rect 13995 10364 14059 10368
rect 13995 10308 13999 10364
rect 13999 10308 14055 10364
rect 14055 10308 14059 10364
rect 13995 10304 14059 10308
rect 6073 9820 6137 9824
rect 6073 9764 6077 9820
rect 6077 9764 6133 9820
rect 6133 9764 6137 9820
rect 6073 9760 6137 9764
rect 6153 9820 6217 9824
rect 6153 9764 6157 9820
rect 6157 9764 6213 9820
rect 6213 9764 6217 9820
rect 6153 9760 6217 9764
rect 6233 9820 6297 9824
rect 6233 9764 6237 9820
rect 6237 9764 6293 9820
rect 6293 9764 6297 9820
rect 6233 9760 6297 9764
rect 6313 9820 6377 9824
rect 6313 9764 6317 9820
rect 6317 9764 6373 9820
rect 6373 9764 6377 9820
rect 6313 9760 6377 9764
rect 11194 9820 11258 9824
rect 11194 9764 11198 9820
rect 11198 9764 11254 9820
rect 11254 9764 11258 9820
rect 11194 9760 11258 9764
rect 11274 9820 11338 9824
rect 11274 9764 11278 9820
rect 11278 9764 11334 9820
rect 11334 9764 11338 9820
rect 11274 9760 11338 9764
rect 11354 9820 11418 9824
rect 11354 9764 11358 9820
rect 11358 9764 11414 9820
rect 11414 9764 11418 9820
rect 11354 9760 11418 9764
rect 11434 9820 11498 9824
rect 11434 9764 11438 9820
rect 11438 9764 11494 9820
rect 11494 9764 11498 9820
rect 11434 9760 11498 9764
rect 3512 9276 3576 9280
rect 3512 9220 3516 9276
rect 3516 9220 3572 9276
rect 3572 9220 3576 9276
rect 3512 9216 3576 9220
rect 3592 9276 3656 9280
rect 3592 9220 3596 9276
rect 3596 9220 3652 9276
rect 3652 9220 3656 9276
rect 3592 9216 3656 9220
rect 3672 9276 3736 9280
rect 3672 9220 3676 9276
rect 3676 9220 3732 9276
rect 3732 9220 3736 9276
rect 3672 9216 3736 9220
rect 3752 9276 3816 9280
rect 3752 9220 3756 9276
rect 3756 9220 3812 9276
rect 3812 9220 3816 9276
rect 3752 9216 3816 9220
rect 8634 9276 8698 9280
rect 8634 9220 8638 9276
rect 8638 9220 8694 9276
rect 8694 9220 8698 9276
rect 8634 9216 8698 9220
rect 8714 9276 8778 9280
rect 8714 9220 8718 9276
rect 8718 9220 8774 9276
rect 8774 9220 8778 9276
rect 8714 9216 8778 9220
rect 8794 9276 8858 9280
rect 8794 9220 8798 9276
rect 8798 9220 8854 9276
rect 8854 9220 8858 9276
rect 8794 9216 8858 9220
rect 8874 9276 8938 9280
rect 8874 9220 8878 9276
rect 8878 9220 8934 9276
rect 8934 9220 8938 9276
rect 8874 9216 8938 9220
rect 13755 9276 13819 9280
rect 13755 9220 13759 9276
rect 13759 9220 13815 9276
rect 13815 9220 13819 9276
rect 13755 9216 13819 9220
rect 13835 9276 13899 9280
rect 13835 9220 13839 9276
rect 13839 9220 13895 9276
rect 13895 9220 13899 9276
rect 13835 9216 13899 9220
rect 13915 9276 13979 9280
rect 13915 9220 13919 9276
rect 13919 9220 13975 9276
rect 13975 9220 13979 9276
rect 13915 9216 13979 9220
rect 13995 9276 14059 9280
rect 13995 9220 13999 9276
rect 13999 9220 14055 9276
rect 14055 9220 14059 9276
rect 13995 9216 14059 9220
rect 6073 8732 6137 8736
rect 6073 8676 6077 8732
rect 6077 8676 6133 8732
rect 6133 8676 6137 8732
rect 6073 8672 6137 8676
rect 6153 8732 6217 8736
rect 6153 8676 6157 8732
rect 6157 8676 6213 8732
rect 6213 8676 6217 8732
rect 6153 8672 6217 8676
rect 6233 8732 6297 8736
rect 6233 8676 6237 8732
rect 6237 8676 6293 8732
rect 6293 8676 6297 8732
rect 6233 8672 6297 8676
rect 6313 8732 6377 8736
rect 6313 8676 6317 8732
rect 6317 8676 6373 8732
rect 6373 8676 6377 8732
rect 6313 8672 6377 8676
rect 11194 8732 11258 8736
rect 11194 8676 11198 8732
rect 11198 8676 11254 8732
rect 11254 8676 11258 8732
rect 11194 8672 11258 8676
rect 11274 8732 11338 8736
rect 11274 8676 11278 8732
rect 11278 8676 11334 8732
rect 11334 8676 11338 8732
rect 11274 8672 11338 8676
rect 11354 8732 11418 8736
rect 11354 8676 11358 8732
rect 11358 8676 11414 8732
rect 11414 8676 11418 8732
rect 11354 8672 11418 8676
rect 11434 8732 11498 8736
rect 11434 8676 11438 8732
rect 11438 8676 11494 8732
rect 11494 8676 11498 8732
rect 11434 8672 11498 8676
rect 3512 8188 3576 8192
rect 3512 8132 3516 8188
rect 3516 8132 3572 8188
rect 3572 8132 3576 8188
rect 3512 8128 3576 8132
rect 3592 8188 3656 8192
rect 3592 8132 3596 8188
rect 3596 8132 3652 8188
rect 3652 8132 3656 8188
rect 3592 8128 3656 8132
rect 3672 8188 3736 8192
rect 3672 8132 3676 8188
rect 3676 8132 3732 8188
rect 3732 8132 3736 8188
rect 3672 8128 3736 8132
rect 3752 8188 3816 8192
rect 3752 8132 3756 8188
rect 3756 8132 3812 8188
rect 3812 8132 3816 8188
rect 3752 8128 3816 8132
rect 8634 8188 8698 8192
rect 8634 8132 8638 8188
rect 8638 8132 8694 8188
rect 8694 8132 8698 8188
rect 8634 8128 8698 8132
rect 8714 8188 8778 8192
rect 8714 8132 8718 8188
rect 8718 8132 8774 8188
rect 8774 8132 8778 8188
rect 8714 8128 8778 8132
rect 8794 8188 8858 8192
rect 8794 8132 8798 8188
rect 8798 8132 8854 8188
rect 8854 8132 8858 8188
rect 8794 8128 8858 8132
rect 8874 8188 8938 8192
rect 8874 8132 8878 8188
rect 8878 8132 8934 8188
rect 8934 8132 8938 8188
rect 8874 8128 8938 8132
rect 13755 8188 13819 8192
rect 13755 8132 13759 8188
rect 13759 8132 13815 8188
rect 13815 8132 13819 8188
rect 13755 8128 13819 8132
rect 13835 8188 13899 8192
rect 13835 8132 13839 8188
rect 13839 8132 13895 8188
rect 13895 8132 13899 8188
rect 13835 8128 13899 8132
rect 13915 8188 13979 8192
rect 13915 8132 13919 8188
rect 13919 8132 13975 8188
rect 13975 8132 13979 8188
rect 13915 8128 13979 8132
rect 13995 8188 14059 8192
rect 13995 8132 13999 8188
rect 13999 8132 14055 8188
rect 14055 8132 14059 8188
rect 13995 8128 14059 8132
rect 6073 7644 6137 7648
rect 6073 7588 6077 7644
rect 6077 7588 6133 7644
rect 6133 7588 6137 7644
rect 6073 7584 6137 7588
rect 6153 7644 6217 7648
rect 6153 7588 6157 7644
rect 6157 7588 6213 7644
rect 6213 7588 6217 7644
rect 6153 7584 6217 7588
rect 6233 7644 6297 7648
rect 6233 7588 6237 7644
rect 6237 7588 6293 7644
rect 6293 7588 6297 7644
rect 6233 7584 6297 7588
rect 6313 7644 6377 7648
rect 6313 7588 6317 7644
rect 6317 7588 6373 7644
rect 6373 7588 6377 7644
rect 6313 7584 6377 7588
rect 11194 7644 11258 7648
rect 11194 7588 11198 7644
rect 11198 7588 11254 7644
rect 11254 7588 11258 7644
rect 11194 7584 11258 7588
rect 11274 7644 11338 7648
rect 11274 7588 11278 7644
rect 11278 7588 11334 7644
rect 11334 7588 11338 7644
rect 11274 7584 11338 7588
rect 11354 7644 11418 7648
rect 11354 7588 11358 7644
rect 11358 7588 11414 7644
rect 11414 7588 11418 7644
rect 11354 7584 11418 7588
rect 11434 7644 11498 7648
rect 11434 7588 11438 7644
rect 11438 7588 11494 7644
rect 11494 7588 11498 7644
rect 11434 7584 11498 7588
rect 3512 7100 3576 7104
rect 3512 7044 3516 7100
rect 3516 7044 3572 7100
rect 3572 7044 3576 7100
rect 3512 7040 3576 7044
rect 3592 7100 3656 7104
rect 3592 7044 3596 7100
rect 3596 7044 3652 7100
rect 3652 7044 3656 7100
rect 3592 7040 3656 7044
rect 3672 7100 3736 7104
rect 3672 7044 3676 7100
rect 3676 7044 3732 7100
rect 3732 7044 3736 7100
rect 3672 7040 3736 7044
rect 3752 7100 3816 7104
rect 3752 7044 3756 7100
rect 3756 7044 3812 7100
rect 3812 7044 3816 7100
rect 3752 7040 3816 7044
rect 8634 7100 8698 7104
rect 8634 7044 8638 7100
rect 8638 7044 8694 7100
rect 8694 7044 8698 7100
rect 8634 7040 8698 7044
rect 8714 7100 8778 7104
rect 8714 7044 8718 7100
rect 8718 7044 8774 7100
rect 8774 7044 8778 7100
rect 8714 7040 8778 7044
rect 8794 7100 8858 7104
rect 8794 7044 8798 7100
rect 8798 7044 8854 7100
rect 8854 7044 8858 7100
rect 8794 7040 8858 7044
rect 8874 7100 8938 7104
rect 8874 7044 8878 7100
rect 8878 7044 8934 7100
rect 8934 7044 8938 7100
rect 8874 7040 8938 7044
rect 13755 7100 13819 7104
rect 13755 7044 13759 7100
rect 13759 7044 13815 7100
rect 13815 7044 13819 7100
rect 13755 7040 13819 7044
rect 13835 7100 13899 7104
rect 13835 7044 13839 7100
rect 13839 7044 13895 7100
rect 13895 7044 13899 7100
rect 13835 7040 13899 7044
rect 13915 7100 13979 7104
rect 13915 7044 13919 7100
rect 13919 7044 13975 7100
rect 13975 7044 13979 7100
rect 13915 7040 13979 7044
rect 13995 7100 14059 7104
rect 13995 7044 13999 7100
rect 13999 7044 14055 7100
rect 14055 7044 14059 7100
rect 13995 7040 14059 7044
rect 6073 6556 6137 6560
rect 6073 6500 6077 6556
rect 6077 6500 6133 6556
rect 6133 6500 6137 6556
rect 6073 6496 6137 6500
rect 6153 6556 6217 6560
rect 6153 6500 6157 6556
rect 6157 6500 6213 6556
rect 6213 6500 6217 6556
rect 6153 6496 6217 6500
rect 6233 6556 6297 6560
rect 6233 6500 6237 6556
rect 6237 6500 6293 6556
rect 6293 6500 6297 6556
rect 6233 6496 6297 6500
rect 6313 6556 6377 6560
rect 6313 6500 6317 6556
rect 6317 6500 6373 6556
rect 6373 6500 6377 6556
rect 6313 6496 6377 6500
rect 11194 6556 11258 6560
rect 11194 6500 11198 6556
rect 11198 6500 11254 6556
rect 11254 6500 11258 6556
rect 11194 6496 11258 6500
rect 11274 6556 11338 6560
rect 11274 6500 11278 6556
rect 11278 6500 11334 6556
rect 11334 6500 11338 6556
rect 11274 6496 11338 6500
rect 11354 6556 11418 6560
rect 11354 6500 11358 6556
rect 11358 6500 11414 6556
rect 11414 6500 11418 6556
rect 11354 6496 11418 6500
rect 11434 6556 11498 6560
rect 11434 6500 11438 6556
rect 11438 6500 11494 6556
rect 11494 6500 11498 6556
rect 11434 6496 11498 6500
rect 8156 6428 8220 6492
rect 3512 6012 3576 6016
rect 3512 5956 3516 6012
rect 3516 5956 3572 6012
rect 3572 5956 3576 6012
rect 3512 5952 3576 5956
rect 3592 6012 3656 6016
rect 3592 5956 3596 6012
rect 3596 5956 3652 6012
rect 3652 5956 3656 6012
rect 3592 5952 3656 5956
rect 3672 6012 3736 6016
rect 3672 5956 3676 6012
rect 3676 5956 3732 6012
rect 3732 5956 3736 6012
rect 3672 5952 3736 5956
rect 3752 6012 3816 6016
rect 3752 5956 3756 6012
rect 3756 5956 3812 6012
rect 3812 5956 3816 6012
rect 3752 5952 3816 5956
rect 8634 6012 8698 6016
rect 8634 5956 8638 6012
rect 8638 5956 8694 6012
rect 8694 5956 8698 6012
rect 8634 5952 8698 5956
rect 8714 6012 8778 6016
rect 8714 5956 8718 6012
rect 8718 5956 8774 6012
rect 8774 5956 8778 6012
rect 8714 5952 8778 5956
rect 8794 6012 8858 6016
rect 8794 5956 8798 6012
rect 8798 5956 8854 6012
rect 8854 5956 8858 6012
rect 8794 5952 8858 5956
rect 8874 6012 8938 6016
rect 8874 5956 8878 6012
rect 8878 5956 8934 6012
rect 8934 5956 8938 6012
rect 8874 5952 8938 5956
rect 13755 6012 13819 6016
rect 13755 5956 13759 6012
rect 13759 5956 13815 6012
rect 13815 5956 13819 6012
rect 13755 5952 13819 5956
rect 13835 6012 13899 6016
rect 13835 5956 13839 6012
rect 13839 5956 13895 6012
rect 13895 5956 13899 6012
rect 13835 5952 13899 5956
rect 13915 6012 13979 6016
rect 13915 5956 13919 6012
rect 13919 5956 13975 6012
rect 13975 5956 13979 6012
rect 13915 5952 13979 5956
rect 13995 6012 14059 6016
rect 13995 5956 13999 6012
rect 13999 5956 14055 6012
rect 14055 5956 14059 6012
rect 13995 5952 14059 5956
rect 6073 5468 6137 5472
rect 6073 5412 6077 5468
rect 6077 5412 6133 5468
rect 6133 5412 6137 5468
rect 6073 5408 6137 5412
rect 6153 5468 6217 5472
rect 6153 5412 6157 5468
rect 6157 5412 6213 5468
rect 6213 5412 6217 5468
rect 6153 5408 6217 5412
rect 6233 5468 6297 5472
rect 6233 5412 6237 5468
rect 6237 5412 6293 5468
rect 6293 5412 6297 5468
rect 6233 5408 6297 5412
rect 6313 5468 6377 5472
rect 6313 5412 6317 5468
rect 6317 5412 6373 5468
rect 6373 5412 6377 5468
rect 6313 5408 6377 5412
rect 11194 5468 11258 5472
rect 11194 5412 11198 5468
rect 11198 5412 11254 5468
rect 11254 5412 11258 5468
rect 11194 5408 11258 5412
rect 11274 5468 11338 5472
rect 11274 5412 11278 5468
rect 11278 5412 11334 5468
rect 11334 5412 11338 5468
rect 11274 5408 11338 5412
rect 11354 5468 11418 5472
rect 11354 5412 11358 5468
rect 11358 5412 11414 5468
rect 11414 5412 11418 5468
rect 11354 5408 11418 5412
rect 11434 5468 11498 5472
rect 11434 5412 11438 5468
rect 11438 5412 11494 5468
rect 11494 5412 11498 5468
rect 11434 5408 11498 5412
rect 3512 4924 3576 4928
rect 3512 4868 3516 4924
rect 3516 4868 3572 4924
rect 3572 4868 3576 4924
rect 3512 4864 3576 4868
rect 3592 4924 3656 4928
rect 3592 4868 3596 4924
rect 3596 4868 3652 4924
rect 3652 4868 3656 4924
rect 3592 4864 3656 4868
rect 3672 4924 3736 4928
rect 3672 4868 3676 4924
rect 3676 4868 3732 4924
rect 3732 4868 3736 4924
rect 3672 4864 3736 4868
rect 3752 4924 3816 4928
rect 3752 4868 3756 4924
rect 3756 4868 3812 4924
rect 3812 4868 3816 4924
rect 3752 4864 3816 4868
rect 8634 4924 8698 4928
rect 8634 4868 8638 4924
rect 8638 4868 8694 4924
rect 8694 4868 8698 4924
rect 8634 4864 8698 4868
rect 8714 4924 8778 4928
rect 8714 4868 8718 4924
rect 8718 4868 8774 4924
rect 8774 4868 8778 4924
rect 8714 4864 8778 4868
rect 8794 4924 8858 4928
rect 8794 4868 8798 4924
rect 8798 4868 8854 4924
rect 8854 4868 8858 4924
rect 8794 4864 8858 4868
rect 8874 4924 8938 4928
rect 8874 4868 8878 4924
rect 8878 4868 8934 4924
rect 8934 4868 8938 4924
rect 8874 4864 8938 4868
rect 13755 4924 13819 4928
rect 13755 4868 13759 4924
rect 13759 4868 13815 4924
rect 13815 4868 13819 4924
rect 13755 4864 13819 4868
rect 13835 4924 13899 4928
rect 13835 4868 13839 4924
rect 13839 4868 13895 4924
rect 13895 4868 13899 4924
rect 13835 4864 13899 4868
rect 13915 4924 13979 4928
rect 13915 4868 13919 4924
rect 13919 4868 13975 4924
rect 13975 4868 13979 4924
rect 13915 4864 13979 4868
rect 13995 4924 14059 4928
rect 13995 4868 13999 4924
rect 13999 4868 14055 4924
rect 14055 4868 14059 4924
rect 13995 4864 14059 4868
rect 6073 4380 6137 4384
rect 6073 4324 6077 4380
rect 6077 4324 6133 4380
rect 6133 4324 6137 4380
rect 6073 4320 6137 4324
rect 6153 4380 6217 4384
rect 6153 4324 6157 4380
rect 6157 4324 6213 4380
rect 6213 4324 6217 4380
rect 6153 4320 6217 4324
rect 6233 4380 6297 4384
rect 6233 4324 6237 4380
rect 6237 4324 6293 4380
rect 6293 4324 6297 4380
rect 6233 4320 6297 4324
rect 6313 4380 6377 4384
rect 6313 4324 6317 4380
rect 6317 4324 6373 4380
rect 6373 4324 6377 4380
rect 6313 4320 6377 4324
rect 11194 4380 11258 4384
rect 11194 4324 11198 4380
rect 11198 4324 11254 4380
rect 11254 4324 11258 4380
rect 11194 4320 11258 4324
rect 11274 4380 11338 4384
rect 11274 4324 11278 4380
rect 11278 4324 11334 4380
rect 11334 4324 11338 4380
rect 11274 4320 11338 4324
rect 11354 4380 11418 4384
rect 11354 4324 11358 4380
rect 11358 4324 11414 4380
rect 11414 4324 11418 4380
rect 11354 4320 11418 4324
rect 11434 4380 11498 4384
rect 11434 4324 11438 4380
rect 11438 4324 11494 4380
rect 11494 4324 11498 4380
rect 11434 4320 11498 4324
rect 3512 3836 3576 3840
rect 3512 3780 3516 3836
rect 3516 3780 3572 3836
rect 3572 3780 3576 3836
rect 3512 3776 3576 3780
rect 3592 3836 3656 3840
rect 3592 3780 3596 3836
rect 3596 3780 3652 3836
rect 3652 3780 3656 3836
rect 3592 3776 3656 3780
rect 3672 3836 3736 3840
rect 3672 3780 3676 3836
rect 3676 3780 3732 3836
rect 3732 3780 3736 3836
rect 3672 3776 3736 3780
rect 3752 3836 3816 3840
rect 3752 3780 3756 3836
rect 3756 3780 3812 3836
rect 3812 3780 3816 3836
rect 3752 3776 3816 3780
rect 8634 3836 8698 3840
rect 8634 3780 8638 3836
rect 8638 3780 8694 3836
rect 8694 3780 8698 3836
rect 8634 3776 8698 3780
rect 8714 3836 8778 3840
rect 8714 3780 8718 3836
rect 8718 3780 8774 3836
rect 8774 3780 8778 3836
rect 8714 3776 8778 3780
rect 8794 3836 8858 3840
rect 8794 3780 8798 3836
rect 8798 3780 8854 3836
rect 8854 3780 8858 3836
rect 8794 3776 8858 3780
rect 8874 3836 8938 3840
rect 8874 3780 8878 3836
rect 8878 3780 8934 3836
rect 8934 3780 8938 3836
rect 8874 3776 8938 3780
rect 13755 3836 13819 3840
rect 13755 3780 13759 3836
rect 13759 3780 13815 3836
rect 13815 3780 13819 3836
rect 13755 3776 13819 3780
rect 13835 3836 13899 3840
rect 13835 3780 13839 3836
rect 13839 3780 13895 3836
rect 13895 3780 13899 3836
rect 13835 3776 13899 3780
rect 13915 3836 13979 3840
rect 13915 3780 13919 3836
rect 13919 3780 13975 3836
rect 13975 3780 13979 3836
rect 13915 3776 13979 3780
rect 13995 3836 14059 3840
rect 13995 3780 13999 3836
rect 13999 3780 14055 3836
rect 14055 3780 14059 3836
rect 13995 3776 14059 3780
rect 6073 3292 6137 3296
rect 6073 3236 6077 3292
rect 6077 3236 6133 3292
rect 6133 3236 6137 3292
rect 6073 3232 6137 3236
rect 6153 3292 6217 3296
rect 6153 3236 6157 3292
rect 6157 3236 6213 3292
rect 6213 3236 6217 3292
rect 6153 3232 6217 3236
rect 6233 3292 6297 3296
rect 6233 3236 6237 3292
rect 6237 3236 6293 3292
rect 6293 3236 6297 3292
rect 6233 3232 6297 3236
rect 6313 3292 6377 3296
rect 6313 3236 6317 3292
rect 6317 3236 6373 3292
rect 6373 3236 6377 3292
rect 6313 3232 6377 3236
rect 11194 3292 11258 3296
rect 11194 3236 11198 3292
rect 11198 3236 11254 3292
rect 11254 3236 11258 3292
rect 11194 3232 11258 3236
rect 11274 3292 11338 3296
rect 11274 3236 11278 3292
rect 11278 3236 11334 3292
rect 11334 3236 11338 3292
rect 11274 3232 11338 3236
rect 11354 3292 11418 3296
rect 11354 3236 11358 3292
rect 11358 3236 11414 3292
rect 11414 3236 11418 3292
rect 11354 3232 11418 3236
rect 11434 3292 11498 3296
rect 11434 3236 11438 3292
rect 11438 3236 11494 3292
rect 11494 3236 11498 3292
rect 11434 3232 11498 3236
rect 8156 2892 8220 2956
rect 3512 2748 3576 2752
rect 3512 2692 3516 2748
rect 3516 2692 3572 2748
rect 3572 2692 3576 2748
rect 3512 2688 3576 2692
rect 3592 2748 3656 2752
rect 3592 2692 3596 2748
rect 3596 2692 3652 2748
rect 3652 2692 3656 2748
rect 3592 2688 3656 2692
rect 3672 2748 3736 2752
rect 3672 2692 3676 2748
rect 3676 2692 3732 2748
rect 3732 2692 3736 2748
rect 3672 2688 3736 2692
rect 3752 2748 3816 2752
rect 3752 2692 3756 2748
rect 3756 2692 3812 2748
rect 3812 2692 3816 2748
rect 3752 2688 3816 2692
rect 8634 2748 8698 2752
rect 8634 2692 8638 2748
rect 8638 2692 8694 2748
rect 8694 2692 8698 2748
rect 8634 2688 8698 2692
rect 8714 2748 8778 2752
rect 8714 2692 8718 2748
rect 8718 2692 8774 2748
rect 8774 2692 8778 2748
rect 8714 2688 8778 2692
rect 8794 2748 8858 2752
rect 8794 2692 8798 2748
rect 8798 2692 8854 2748
rect 8854 2692 8858 2748
rect 8794 2688 8858 2692
rect 8874 2748 8938 2752
rect 8874 2692 8878 2748
rect 8878 2692 8934 2748
rect 8934 2692 8938 2748
rect 8874 2688 8938 2692
rect 13755 2748 13819 2752
rect 13755 2692 13759 2748
rect 13759 2692 13815 2748
rect 13815 2692 13819 2748
rect 13755 2688 13819 2692
rect 13835 2748 13899 2752
rect 13835 2692 13839 2748
rect 13839 2692 13895 2748
rect 13895 2692 13899 2748
rect 13835 2688 13899 2692
rect 13915 2748 13979 2752
rect 13915 2692 13919 2748
rect 13919 2692 13975 2748
rect 13975 2692 13979 2748
rect 13915 2688 13979 2692
rect 13995 2748 14059 2752
rect 13995 2692 13999 2748
rect 13999 2692 14055 2748
rect 14055 2692 14059 2748
rect 13995 2688 14059 2692
rect 6073 2204 6137 2208
rect 6073 2148 6077 2204
rect 6077 2148 6133 2204
rect 6133 2148 6137 2204
rect 6073 2144 6137 2148
rect 6153 2204 6217 2208
rect 6153 2148 6157 2204
rect 6157 2148 6213 2204
rect 6213 2148 6217 2204
rect 6153 2144 6217 2148
rect 6233 2204 6297 2208
rect 6233 2148 6237 2204
rect 6237 2148 6293 2204
rect 6293 2148 6297 2204
rect 6233 2144 6297 2148
rect 6313 2204 6377 2208
rect 6313 2148 6317 2204
rect 6317 2148 6373 2204
rect 6373 2148 6377 2204
rect 6313 2144 6377 2148
rect 11194 2204 11258 2208
rect 11194 2148 11198 2204
rect 11198 2148 11254 2204
rect 11254 2148 11258 2204
rect 11194 2144 11258 2148
rect 11274 2204 11338 2208
rect 11274 2148 11278 2204
rect 11278 2148 11334 2204
rect 11334 2148 11338 2204
rect 11274 2144 11338 2148
rect 11354 2204 11418 2208
rect 11354 2148 11358 2204
rect 11358 2148 11414 2204
rect 11414 2148 11418 2204
rect 11354 2144 11418 2148
rect 11434 2204 11498 2208
rect 11434 2148 11438 2204
rect 11438 2148 11494 2204
rect 11494 2148 11498 2204
rect 11434 2144 11498 2148
<< metal4 >>
rect 3504 16896 3824 17456
rect 3504 16832 3512 16896
rect 3576 16832 3592 16896
rect 3656 16832 3672 16896
rect 3736 16832 3752 16896
rect 3816 16832 3824 16896
rect 3504 15808 3824 16832
rect 3504 15744 3512 15808
rect 3576 15744 3592 15808
rect 3656 15744 3672 15808
rect 3736 15744 3752 15808
rect 3816 15744 3824 15808
rect 3504 14939 3824 15744
rect 3504 14720 3546 14939
rect 3782 14720 3824 14939
rect 3504 14656 3512 14720
rect 3576 14656 3592 14703
rect 3656 14656 3672 14703
rect 3736 14656 3752 14703
rect 3816 14656 3824 14720
rect 3504 13632 3824 14656
rect 3504 13568 3512 13632
rect 3576 13568 3592 13632
rect 3656 13568 3672 13632
rect 3736 13568 3752 13632
rect 3816 13568 3824 13632
rect 3504 12544 3824 13568
rect 3504 12480 3512 12544
rect 3576 12480 3592 12544
rect 3656 12480 3672 12544
rect 3736 12480 3752 12544
rect 3816 12480 3824 12544
rect 3504 11456 3824 12480
rect 3504 11392 3512 11456
rect 3576 11392 3592 11456
rect 3656 11392 3672 11456
rect 3736 11392 3752 11456
rect 3816 11392 3824 11456
rect 3504 10368 3824 11392
rect 3504 10304 3512 10368
rect 3576 10304 3592 10368
rect 3656 10304 3672 10368
rect 3736 10304 3752 10368
rect 3816 10304 3824 10368
rect 3504 9862 3824 10304
rect 3504 9626 3546 9862
rect 3782 9626 3824 9862
rect 3504 9280 3824 9626
rect 3504 9216 3512 9280
rect 3576 9216 3592 9280
rect 3656 9216 3672 9280
rect 3736 9216 3752 9280
rect 3816 9216 3824 9280
rect 3504 8192 3824 9216
rect 3504 8128 3512 8192
rect 3576 8128 3592 8192
rect 3656 8128 3672 8192
rect 3736 8128 3752 8192
rect 3816 8128 3824 8192
rect 3504 7104 3824 8128
rect 3504 7040 3512 7104
rect 3576 7040 3592 7104
rect 3656 7040 3672 7104
rect 3736 7040 3752 7104
rect 3816 7040 3824 7104
rect 3504 6016 3824 7040
rect 3504 5952 3512 6016
rect 3576 5952 3592 6016
rect 3656 5952 3672 6016
rect 3736 5952 3752 6016
rect 3816 5952 3824 6016
rect 3504 4928 3824 5952
rect 3504 4864 3512 4928
rect 3576 4864 3592 4928
rect 3656 4864 3672 4928
rect 3736 4864 3752 4928
rect 3816 4864 3824 4928
rect 3504 4784 3824 4864
rect 3504 4548 3546 4784
rect 3782 4548 3824 4784
rect 3504 3840 3824 4548
rect 3504 3776 3512 3840
rect 3576 3776 3592 3840
rect 3656 3776 3672 3840
rect 3736 3776 3752 3840
rect 3816 3776 3824 3840
rect 3504 2752 3824 3776
rect 3504 2688 3512 2752
rect 3576 2688 3592 2752
rect 3656 2688 3672 2752
rect 3736 2688 3752 2752
rect 3816 2688 3824 2752
rect 3504 2128 3824 2688
rect 6065 17440 6385 17456
rect 6065 17376 6073 17440
rect 6137 17376 6153 17440
rect 6217 17376 6233 17440
rect 6297 17376 6313 17440
rect 6377 17376 6385 17440
rect 6065 16352 6385 17376
rect 6065 16288 6073 16352
rect 6137 16288 6153 16352
rect 6217 16288 6233 16352
rect 6297 16288 6313 16352
rect 6377 16288 6385 16352
rect 6065 15264 6385 16288
rect 6065 15200 6073 15264
rect 6137 15200 6153 15264
rect 6217 15200 6233 15264
rect 6297 15200 6313 15264
rect 6377 15200 6385 15264
rect 6065 14176 6385 15200
rect 6065 14112 6073 14176
rect 6137 14112 6153 14176
rect 6217 14112 6233 14176
rect 6297 14112 6313 14176
rect 6377 14112 6385 14176
rect 6065 13088 6385 14112
rect 6065 13024 6073 13088
rect 6137 13024 6153 13088
rect 6217 13024 6233 13088
rect 6297 13024 6313 13088
rect 6377 13024 6385 13088
rect 6065 12400 6385 13024
rect 6065 12164 6107 12400
rect 6343 12164 6385 12400
rect 6065 12000 6385 12164
rect 6065 11936 6073 12000
rect 6137 11936 6153 12000
rect 6217 11936 6233 12000
rect 6297 11936 6313 12000
rect 6377 11936 6385 12000
rect 6065 10912 6385 11936
rect 6065 10848 6073 10912
rect 6137 10848 6153 10912
rect 6217 10848 6233 10912
rect 6297 10848 6313 10912
rect 6377 10848 6385 10912
rect 6065 9824 6385 10848
rect 6065 9760 6073 9824
rect 6137 9760 6153 9824
rect 6217 9760 6233 9824
rect 6297 9760 6313 9824
rect 6377 9760 6385 9824
rect 6065 8736 6385 9760
rect 6065 8672 6073 8736
rect 6137 8672 6153 8736
rect 6217 8672 6233 8736
rect 6297 8672 6313 8736
rect 6377 8672 6385 8736
rect 6065 7648 6385 8672
rect 6065 7584 6073 7648
rect 6137 7584 6153 7648
rect 6217 7584 6233 7648
rect 6297 7584 6313 7648
rect 6377 7584 6385 7648
rect 6065 7323 6385 7584
rect 6065 7087 6107 7323
rect 6343 7087 6385 7323
rect 6065 6560 6385 7087
rect 6065 6496 6073 6560
rect 6137 6496 6153 6560
rect 6217 6496 6233 6560
rect 6297 6496 6313 6560
rect 6377 6496 6385 6560
rect 6065 5472 6385 6496
rect 8626 16896 8946 17456
rect 8626 16832 8634 16896
rect 8698 16832 8714 16896
rect 8778 16832 8794 16896
rect 8858 16832 8874 16896
rect 8938 16832 8946 16896
rect 8626 15808 8946 16832
rect 8626 15744 8634 15808
rect 8698 15744 8714 15808
rect 8778 15744 8794 15808
rect 8858 15744 8874 15808
rect 8938 15744 8946 15808
rect 8626 14939 8946 15744
rect 8626 14720 8668 14939
rect 8904 14720 8946 14939
rect 8626 14656 8634 14720
rect 8698 14656 8714 14703
rect 8778 14656 8794 14703
rect 8858 14656 8874 14703
rect 8938 14656 8946 14720
rect 8626 13632 8946 14656
rect 8626 13568 8634 13632
rect 8698 13568 8714 13632
rect 8778 13568 8794 13632
rect 8858 13568 8874 13632
rect 8938 13568 8946 13632
rect 8626 12544 8946 13568
rect 8626 12480 8634 12544
rect 8698 12480 8714 12544
rect 8778 12480 8794 12544
rect 8858 12480 8874 12544
rect 8938 12480 8946 12544
rect 8626 11456 8946 12480
rect 8626 11392 8634 11456
rect 8698 11392 8714 11456
rect 8778 11392 8794 11456
rect 8858 11392 8874 11456
rect 8938 11392 8946 11456
rect 8626 10368 8946 11392
rect 8626 10304 8634 10368
rect 8698 10304 8714 10368
rect 8778 10304 8794 10368
rect 8858 10304 8874 10368
rect 8938 10304 8946 10368
rect 8626 9862 8946 10304
rect 8626 9626 8668 9862
rect 8904 9626 8946 9862
rect 8626 9280 8946 9626
rect 8626 9216 8634 9280
rect 8698 9216 8714 9280
rect 8778 9216 8794 9280
rect 8858 9216 8874 9280
rect 8938 9216 8946 9280
rect 8626 8192 8946 9216
rect 8626 8128 8634 8192
rect 8698 8128 8714 8192
rect 8778 8128 8794 8192
rect 8858 8128 8874 8192
rect 8938 8128 8946 8192
rect 8626 7104 8946 8128
rect 8626 7040 8634 7104
rect 8698 7040 8714 7104
rect 8778 7040 8794 7104
rect 8858 7040 8874 7104
rect 8938 7040 8946 7104
rect 8155 6492 8221 6493
rect 8155 6428 8156 6492
rect 8220 6428 8221 6492
rect 8155 6427 8221 6428
rect 6065 5408 6073 5472
rect 6137 5408 6153 5472
rect 6217 5408 6233 5472
rect 6297 5408 6313 5472
rect 6377 5408 6385 5472
rect 6065 4384 6385 5408
rect 6065 4320 6073 4384
rect 6137 4320 6153 4384
rect 6217 4320 6233 4384
rect 6297 4320 6313 4384
rect 6377 4320 6385 4384
rect 6065 3296 6385 4320
rect 6065 3232 6073 3296
rect 6137 3232 6153 3296
rect 6217 3232 6233 3296
rect 6297 3232 6313 3296
rect 6377 3232 6385 3296
rect 6065 2208 6385 3232
rect 8158 2957 8218 6427
rect 8626 6016 8946 7040
rect 8626 5952 8634 6016
rect 8698 5952 8714 6016
rect 8778 5952 8794 6016
rect 8858 5952 8874 6016
rect 8938 5952 8946 6016
rect 8626 4928 8946 5952
rect 8626 4864 8634 4928
rect 8698 4864 8714 4928
rect 8778 4864 8794 4928
rect 8858 4864 8874 4928
rect 8938 4864 8946 4928
rect 8626 4784 8946 4864
rect 8626 4548 8668 4784
rect 8904 4548 8946 4784
rect 8626 3840 8946 4548
rect 8626 3776 8634 3840
rect 8698 3776 8714 3840
rect 8778 3776 8794 3840
rect 8858 3776 8874 3840
rect 8938 3776 8946 3840
rect 8155 2956 8221 2957
rect 8155 2892 8156 2956
rect 8220 2892 8221 2956
rect 8155 2891 8221 2892
rect 6065 2144 6073 2208
rect 6137 2144 6153 2208
rect 6217 2144 6233 2208
rect 6297 2144 6313 2208
rect 6377 2144 6385 2208
rect 6065 2128 6385 2144
rect 8626 2752 8946 3776
rect 8626 2688 8634 2752
rect 8698 2688 8714 2752
rect 8778 2688 8794 2752
rect 8858 2688 8874 2752
rect 8938 2688 8946 2752
rect 8626 2128 8946 2688
rect 11186 17440 11506 17456
rect 11186 17376 11194 17440
rect 11258 17376 11274 17440
rect 11338 17376 11354 17440
rect 11418 17376 11434 17440
rect 11498 17376 11506 17440
rect 11186 16352 11506 17376
rect 11186 16288 11194 16352
rect 11258 16288 11274 16352
rect 11338 16288 11354 16352
rect 11418 16288 11434 16352
rect 11498 16288 11506 16352
rect 11186 15264 11506 16288
rect 11186 15200 11194 15264
rect 11258 15200 11274 15264
rect 11338 15200 11354 15264
rect 11418 15200 11434 15264
rect 11498 15200 11506 15264
rect 11186 14176 11506 15200
rect 11186 14112 11194 14176
rect 11258 14112 11274 14176
rect 11338 14112 11354 14176
rect 11418 14112 11434 14176
rect 11498 14112 11506 14176
rect 11186 13088 11506 14112
rect 11186 13024 11194 13088
rect 11258 13024 11274 13088
rect 11338 13024 11354 13088
rect 11418 13024 11434 13088
rect 11498 13024 11506 13088
rect 11186 12400 11506 13024
rect 11186 12164 11228 12400
rect 11464 12164 11506 12400
rect 11186 12000 11506 12164
rect 11186 11936 11194 12000
rect 11258 11936 11274 12000
rect 11338 11936 11354 12000
rect 11418 11936 11434 12000
rect 11498 11936 11506 12000
rect 11186 10912 11506 11936
rect 11186 10848 11194 10912
rect 11258 10848 11274 10912
rect 11338 10848 11354 10912
rect 11418 10848 11434 10912
rect 11498 10848 11506 10912
rect 11186 9824 11506 10848
rect 11186 9760 11194 9824
rect 11258 9760 11274 9824
rect 11338 9760 11354 9824
rect 11418 9760 11434 9824
rect 11498 9760 11506 9824
rect 11186 8736 11506 9760
rect 11186 8672 11194 8736
rect 11258 8672 11274 8736
rect 11338 8672 11354 8736
rect 11418 8672 11434 8736
rect 11498 8672 11506 8736
rect 11186 7648 11506 8672
rect 11186 7584 11194 7648
rect 11258 7584 11274 7648
rect 11338 7584 11354 7648
rect 11418 7584 11434 7648
rect 11498 7584 11506 7648
rect 11186 7323 11506 7584
rect 11186 7087 11228 7323
rect 11464 7087 11506 7323
rect 11186 6560 11506 7087
rect 11186 6496 11194 6560
rect 11258 6496 11274 6560
rect 11338 6496 11354 6560
rect 11418 6496 11434 6560
rect 11498 6496 11506 6560
rect 11186 5472 11506 6496
rect 11186 5408 11194 5472
rect 11258 5408 11274 5472
rect 11338 5408 11354 5472
rect 11418 5408 11434 5472
rect 11498 5408 11506 5472
rect 11186 4384 11506 5408
rect 11186 4320 11194 4384
rect 11258 4320 11274 4384
rect 11338 4320 11354 4384
rect 11418 4320 11434 4384
rect 11498 4320 11506 4384
rect 11186 3296 11506 4320
rect 11186 3232 11194 3296
rect 11258 3232 11274 3296
rect 11338 3232 11354 3296
rect 11418 3232 11434 3296
rect 11498 3232 11506 3296
rect 11186 2208 11506 3232
rect 11186 2144 11194 2208
rect 11258 2144 11274 2208
rect 11338 2144 11354 2208
rect 11418 2144 11434 2208
rect 11498 2144 11506 2208
rect 11186 2128 11506 2144
rect 13747 16896 14067 17456
rect 13747 16832 13755 16896
rect 13819 16832 13835 16896
rect 13899 16832 13915 16896
rect 13979 16832 13995 16896
rect 14059 16832 14067 16896
rect 13747 15808 14067 16832
rect 13747 15744 13755 15808
rect 13819 15744 13835 15808
rect 13899 15744 13915 15808
rect 13979 15744 13995 15808
rect 14059 15744 14067 15808
rect 13747 14939 14067 15744
rect 13747 14720 13789 14939
rect 14025 14720 14067 14939
rect 13747 14656 13755 14720
rect 13819 14656 13835 14703
rect 13899 14656 13915 14703
rect 13979 14656 13995 14703
rect 14059 14656 14067 14720
rect 13747 13632 14067 14656
rect 13747 13568 13755 13632
rect 13819 13568 13835 13632
rect 13899 13568 13915 13632
rect 13979 13568 13995 13632
rect 14059 13568 14067 13632
rect 13747 12544 14067 13568
rect 13747 12480 13755 12544
rect 13819 12480 13835 12544
rect 13899 12480 13915 12544
rect 13979 12480 13995 12544
rect 14059 12480 14067 12544
rect 13747 11456 14067 12480
rect 13747 11392 13755 11456
rect 13819 11392 13835 11456
rect 13899 11392 13915 11456
rect 13979 11392 13995 11456
rect 14059 11392 14067 11456
rect 13747 10368 14067 11392
rect 13747 10304 13755 10368
rect 13819 10304 13835 10368
rect 13899 10304 13915 10368
rect 13979 10304 13995 10368
rect 14059 10304 14067 10368
rect 13747 9862 14067 10304
rect 13747 9626 13789 9862
rect 14025 9626 14067 9862
rect 13747 9280 14067 9626
rect 13747 9216 13755 9280
rect 13819 9216 13835 9280
rect 13899 9216 13915 9280
rect 13979 9216 13995 9280
rect 14059 9216 14067 9280
rect 13747 8192 14067 9216
rect 13747 8128 13755 8192
rect 13819 8128 13835 8192
rect 13899 8128 13915 8192
rect 13979 8128 13995 8192
rect 14059 8128 14067 8192
rect 13747 7104 14067 8128
rect 13747 7040 13755 7104
rect 13819 7040 13835 7104
rect 13899 7040 13915 7104
rect 13979 7040 13995 7104
rect 14059 7040 14067 7104
rect 13747 6016 14067 7040
rect 13747 5952 13755 6016
rect 13819 5952 13835 6016
rect 13899 5952 13915 6016
rect 13979 5952 13995 6016
rect 14059 5952 14067 6016
rect 13747 4928 14067 5952
rect 13747 4864 13755 4928
rect 13819 4864 13835 4928
rect 13899 4864 13915 4928
rect 13979 4864 13995 4928
rect 14059 4864 14067 4928
rect 13747 4784 14067 4864
rect 13747 4548 13789 4784
rect 14025 4548 14067 4784
rect 13747 3840 14067 4548
rect 13747 3776 13755 3840
rect 13819 3776 13835 3840
rect 13899 3776 13915 3840
rect 13979 3776 13995 3840
rect 14059 3776 14067 3840
rect 13747 2752 14067 3776
rect 13747 2688 13755 2752
rect 13819 2688 13835 2752
rect 13899 2688 13915 2752
rect 13979 2688 13995 2752
rect 14059 2688 14067 2752
rect 13747 2128 14067 2688
<< via4 >>
rect 3546 14720 3782 14939
rect 3546 14703 3576 14720
rect 3576 14703 3592 14720
rect 3592 14703 3656 14720
rect 3656 14703 3672 14720
rect 3672 14703 3736 14720
rect 3736 14703 3752 14720
rect 3752 14703 3782 14720
rect 3546 9626 3782 9862
rect 3546 4548 3782 4784
rect 6107 12164 6343 12400
rect 6107 7087 6343 7323
rect 8668 14720 8904 14939
rect 8668 14703 8698 14720
rect 8698 14703 8714 14720
rect 8714 14703 8778 14720
rect 8778 14703 8794 14720
rect 8794 14703 8858 14720
rect 8858 14703 8874 14720
rect 8874 14703 8904 14720
rect 8668 9626 8904 9862
rect 8668 4548 8904 4784
rect 11228 12164 11464 12400
rect 11228 7087 11464 7323
rect 13789 14720 14025 14939
rect 13789 14703 13819 14720
rect 13819 14703 13835 14720
rect 13835 14703 13899 14720
rect 13899 14703 13915 14720
rect 13915 14703 13979 14720
rect 13979 14703 13995 14720
rect 13995 14703 14025 14720
rect 13789 9626 14025 9862
rect 13789 4548 14025 4784
<< metal5 >>
rect 1104 14939 16468 14981
rect 1104 14703 3546 14939
rect 3782 14703 8668 14939
rect 8904 14703 13789 14939
rect 14025 14703 16468 14939
rect 1104 14661 16468 14703
rect 1104 12400 16468 12442
rect 1104 12164 6107 12400
rect 6343 12164 11228 12400
rect 11464 12164 16468 12400
rect 1104 12122 16468 12164
rect 1104 9862 16468 9904
rect 1104 9626 3546 9862
rect 3782 9626 8668 9862
rect 8904 9626 13789 9862
rect 14025 9626 16468 9862
rect 1104 9584 16468 9626
rect 1104 7323 16468 7366
rect 1104 7087 6107 7323
rect 6343 7087 11228 7323
rect 11464 7087 16468 7323
rect 1104 7045 16468 7087
rect 1104 4784 16468 4826
rect 1104 4548 3546 4784
rect 3782 4548 8668 4784
rect 8904 4548 13789 4784
rect 14025 4548 16468 4784
rect 1104 4506 16468 4548
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1629484573
transform 1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1629484573
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1629484573
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _620_
timestamp 1629484573
transform -1 0 2116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1629484573
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1629484573
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21
timestamp 1629484573
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_18
timestamp 1629484573
transform 1 0 2760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _610_
timestamp 1629484573
transform -1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _617_
timestamp 1629484573
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output20
timestamp 1629484573
transform -1 0 3036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1629484573
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1629484573
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37
timestamp 1629484573
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1629484573
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_37
timestamp 1629484573
transform 1 0 4508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1629484573
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _626_
timestamp 1629484573
transform 1 0 3864 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output21
timestamp 1629484573
transform -1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44
timestamp 1629484573
transform 1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_43
timestamp 1629484573
transform 1 0 5060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _588_
timestamp 1629484573
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _614_
timestamp 1629484573
transform 1 0 5152 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output24
timestamp 1629484573
transform -1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1629484573
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64
timestamp 1629484573
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1629484573
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1629484573
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1629484573
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1629484573
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _589_
timestamp 1629484573
transform 1 0 6900 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _621_
timestamp 1629484573
transform -1 0 6992 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71
timestamp 1629484573
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1629484573
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _569_
timestamp 1629484573
transform -1 0 7636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _613_
timestamp 1629484573
transform 1 0 8004 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _622_
timestamp 1629484573
transform 1 0 8004 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1629484573
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_83
timestamp 1629484573
transform 1 0 8740 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1629484573
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _584_
timestamp 1629484573
transform -1 0 9384 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102
timestamp 1629484573
transform 1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1629484573
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1629484573
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_1  _623_
timestamp 1629484573
transform 1 0 9752 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_2  _628_
timestamp 1629484573
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1629484573
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1629484573
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1629484573
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1629484573
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1629484573
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1629484573
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _451_
timestamp 1629484573
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121
timestamp 1629484573
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128
timestamp 1629484573
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_116
timestamp 1629484573
transform 1 0 11776 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _315_
timestamp 1629484573
transform 1 0 12144 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _560_
timestamp 1629484573
transform -1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output29
timestamp 1629484573
transform -1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1629484573
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1629484573
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141
timestamp 1629484573
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1629484573
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1629484573
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1629484573
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _454_
timestamp 1629484573
transform 1 0 13340 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _561_
timestamp 1629484573
transform -1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145
timestamp 1629484573
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152
timestamp 1629484573
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_150
timestamp 1629484573
transform 1 0 14904 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1629484573
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _415_
timestamp 1629484573
transform -1 0 14444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _452_
timestamp 1629484573
transform 1 0 14444 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_0_160
timestamp 1629484573
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_160
timestamp 1629484573
transform 1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1629484573
transform -1 0 16468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1629484573
transform -1 0 16468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output19
timestamp 1629484573
transform -1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output23
timestamp 1629484573
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_6
timestamp 1629484573
transform 1 0 1656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1629484573
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _612_
timestamp 1629484573
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_2  _625_
timestamp 1629484573
transform 1 0 2024 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1629484573
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1629484573
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1629484573
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _624_
timestamp 1629484573
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1629484573
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1629484573
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _585_
timestamp 1629484573
transform -1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _611_
timestamp 1629484573
transform 1 0 5612 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_56
timestamp 1629484573
transform 1 0 6256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _590_
timestamp 1629484573
transform -1 0 7084 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_2_65
timestamp 1629484573
transform 1 0 7084 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _586_
timestamp 1629484573
transform 1 0 7636 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1629484573
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1629484573
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _608_
timestamp 1629484573
transform -1 0 9568 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_2_92
timestamp 1629484573
transform 1 0 9568 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_98
timestamp 1629484573
transform 1 0 10120 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _564_
timestamp 1629484573
transform -1 0 10764 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_105
timestamp 1629484573
transform 1 0 10764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _562_
timestamp 1629484573
transform 1 0 11132 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_116
timestamp 1629484573
transform 1 0 11776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_120
timestamp 1629484573
transform 1 0 12144 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_124
timestamp 1629484573
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1629484573
transform -1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _487_
timestamp 1629484573
transform 1 0 12880 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1629484573
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1629484573
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1629484573
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_1  _453_
timestamp 1629484573
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1629484573
transform 1 0 14812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1629484573
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_156
timestamp 1629484573
transform 1 0 15456 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1629484573
transform -1 0 16468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_10
timestamp 1629484573
transform 1 0 2024 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1629484573
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1629484573
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _619_
timestamp 1629484573
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_18
timestamp 1629484573
transform 1 0 2760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_22
timestamp 1629484573
transform 1 0 3128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _599_
timestamp 1629484573
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_29
timestamp 1629484573
transform 1 0 3772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1629484573
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _587_
timestamp 1629484573
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _591_
timestamp 1629484573
transform -1 0 3772 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_43
timestamp 1629484573
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1629484573
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _573_
timestamp 1629484573
transform -1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _592_
timestamp 1629484573
transform 1 0 5428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1629484573
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57
timestamp 1629484573
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1629484573
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _545_
timestamp 1629484573
transform -1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_66
timestamp 1629484573
transform 1 0 7176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _469_
timestamp 1629484573
transform 1 0 7544 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_3_80
timestamp 1629484573
transform 1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _609_
timestamp 1629484573
transform 1 0 8832 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_3_101
timestamp 1629484573
transform 1 0 10396 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_91
timestamp 1629484573
transform 1 0 9476 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _627_
timestamp 1629484573
transform -1 0 10396 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1629484573
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1629484573
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1629484573
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _563_
timestamp 1629484573
transform -1 0 12052 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_119
timestamp 1629484573
transform 1 0 12052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_126
timestamp 1629484573
transform 1 0 12696 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1629484573
transform -1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_130
timestamp 1629484573
transform 1 0 13064 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_134
timestamp 1629484573
transform 1 0 13432 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1629484573
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp 1629484573
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _418_
timestamp 1629484573
transform 1 0 14996 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _448_
timestamp 1629484573
transform -1 0 14628 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_3_156
timestamp 1629484573
transform 1 0 15456 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1629484573
transform -1 0 16468 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1629484573
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1629484573
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _607_
timestamp 1629484573
transform -1 0 2300 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_4_13
timestamp 1629484573
transform 1 0 2300 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1629484573
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _593_
timestamp 1629484573
transform -1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_36
timestamp 1629484573
transform 1 0 4416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1629484573
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _600_
timestamp 1629484573
transform 1 0 3772 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_4_47
timestamp 1629484573
transform 1 0 5428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _572_
timestamp 1629484573
transform -1 0 6256 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _615_
timestamp 1629484573
transform 1 0 4784 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_4_56
timestamp 1629484573
transform 1 0 6256 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_64
timestamp 1629484573
transform 1 0 6992 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_69
timestamp 1629484573
transform 1 0 7452 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1629484573
transform 1 0 7176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _543_
timestamp 1629484573
transform -1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1629484573
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1629484573
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _404_
timestamp 1629484573
transform 1 0 8924 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_4_95
timestamp 1629484573
transform 1 0 9844 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _514_
timestamp 1629484573
transform -1 0 10856 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_4_106
timestamp 1629484573
transform 1 0 10856 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _541_
timestamp 1629484573
transform 1 0 11224 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1629484573
transform 1 0 11868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_125
timestamp 1629484573
transform 1 0 12604 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _347_
timestamp 1629484573
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1629484573
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1629484573
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _311_
timestamp 1629484573
transform -1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _519_
timestamp 1629484573
transform -1 0 13616 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1629484573
transform 1 0 14352 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_148
timestamp 1629484573
transform 1 0 14720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _378_
timestamp 1629484573
transform 1 0 14812 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_4_159
timestamp 1629484573
transform 1 0 15732 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_163
timestamp 1629484573
transform 1 0 16100 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1629484573
transform -1 0 16468 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1629484573
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1629484573
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1629484573
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _601_
timestamp 1629484573
transform -1 0 2392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _606_
timestamp 1629484573
transform -1 0 1748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_14
timestamp 1629484573
transform 1 0 2392 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_20
timestamp 1629484573
transform 1 0 2944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _598_
timestamp 1629484573
transform -1 0 3496 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_5_26
timestamp 1629484573
transform 1 0 3496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1629484573
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _596_
timestamp 1629484573
transform 1 0 3864 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1629484573
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _594_
timestamp 1629484573
transform -1 0 5612 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1629484573
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1629484573
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1629484573
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _595_
timestamp 1629484573
transform 1 0 6716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 1629484573
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_76
timestamp 1629484573
transform 1 0 8096 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _435_
timestamp 1629484573
transform 1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _544_
timestamp 1629484573
transform 1 0 8648 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_5_92
timestamp 1629484573
transform 1 0 9568 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_98
timestamp 1629484573
transform 1 0 10120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__and4_1  _542_
timestamp 1629484573
transform 1 0 10212 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1629484573
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1629484573
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1629484573
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _512_
timestamp 1629484573
transform 1 0 11592 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_5_121
timestamp 1629484573
transform 1 0 12236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_127
timestamp 1629484573
transform 1 0 12788 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _484_
timestamp 1629484573
transform 1 0 12880 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1629484573
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _417_
timestamp 1629484573
transform 1 0 13892 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_5_146
timestamp 1629484573
transform 1 0 14536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _324_
timestamp 1629484573
transform 1 0 14904 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_5_160
timestamp 1629484573
transform 1 0 15824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1629484573
transform -1 0 16468 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_6
timestamp 1629484573
transform 1 0 1656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1629484573
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1629484573
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _616_
timestamp 1629484573
transform -1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _618_
timestamp 1629484573
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1629484573
transform 1 0 1380 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1629484573
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1629484573
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_13
timestamp 1629484573
transform 1 0 2300 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_21
timestamp 1629484573
transform 1 0 3036 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_1  _576_
timestamp 1629484573
transform 1 0 3220 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _597_
timestamp 1629484573
transform 1 0 2668 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1629484573
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_31
timestamp 1629484573
transform 1 0 3956 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1629484573
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _575_
timestamp 1629484573
transform 1 0 4324 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp 1629484573
transform 1 0 4968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_39
timestamp 1629484573
transform 1 0 4692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_49
timestamp 1629484573
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _548_
timestamp 1629484573
transform 1 0 4876 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _574_
timestamp 1629484573
transform 1 0 5336 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_52
timestamp 1629484573
transform 1 0 5888 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1629484573
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_60
timestamp 1629484573
transform 1 0 6624 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1629484573
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _566_
timestamp 1629484573
transform -1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _570_
timestamp 1629484573
transform -1 0 7452 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _571_
timestamp 1629484573
transform 1 0 6624 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_68
timestamp 1629484573
transform 1 0 7360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_69
timestamp 1629484573
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _536_
timestamp 1629484573
transform -1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _568_
timestamp 1629484573
transform -1 0 8464 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1629484573
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1629484573
transform 1 0 8280 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_85
timestamp 1629484573
transform 1 0 8924 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1629484573
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _515_
timestamp 1629484573
transform -1 0 9568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _535_
timestamp 1629484573
transform -1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _546_
timestamp 1629484573
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_93
timestamp 1629484573
transform 1 0 9660 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_92
timestamp 1629484573
transform 1 0 9568 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _513_
timestamp 1629484573
transform 1 0 10212 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _534_
timestamp 1629484573
transform 1 0 9936 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_106
timestamp 1629484573
transform 1 0 10856 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_103
timestamp 1629484573
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1629484573
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_113
timestamp 1629484573
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1629484573
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _565_
timestamp 1629484573
transform 1 0 11224 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_6_117
timestamp 1629484573
transform 1 0 11868 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_125
timestamp 1629484573
transform 1 0 12604 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_124
timestamp 1629484573
transform 1 0 12512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _485_
timestamp 1629484573
transform -1 0 13432 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _486_
timestamp 1629484573
transform -1 0 12512 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _547_
timestamp 1629484573
transform 1 0 12880 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 1629484573
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1629484573
transform 1 0 13616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1629484573
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _447_
timestamp 1629484573
transform -1 0 14536 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  output32
timestamp 1629484573
transform 1 0 13984 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 1629484573
transform 1 0 14536 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_144
timestamp 1629484573
transform 1 0 14352 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _416_
timestamp 1629484573
transform -1 0 15548 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _455_
timestamp 1629484573
transform 1 0 14720 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_157
timestamp 1629484573
transform 1 0 15548 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_163
timestamp 1629484573
transform 1 0 16100 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_156
timestamp 1629484573
transform 1 0 15456 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1629484573
transform -1 0 16468 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1629484573
transform -1 0 16468 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_6
timestamp 1629484573
transform 1 0 1656 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1629484573
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1629484573
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1629484573
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _577_
timestamp 1629484573
transform 1 0 2392 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_37
timestamp 1629484573
transform 1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1629484573
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _549_
timestamp 1629484573
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_45
timestamp 1629484573
transform 1 0 5244 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_49
timestamp 1629484573
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _567_
timestamp 1629484573
transform -1 0 5612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_56
timestamp 1629484573
transform 1 0 6256 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _538_
timestamp 1629484573
transform -1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _559_
timestamp 1629484573
transform 1 0 6624 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_68
timestamp 1629484573
transform 1 0 7360 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _537_
timestamp 1629484573
transform 1 0 7728 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1629484573
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1629484573
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1629484573
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _516_
timestamp 1629484573
transform -1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_92
timestamp 1629484573
transform 1 0 9568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _386_
timestamp 1629484573
transform 1 0 9936 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_8_106
timestamp 1629484573
transform 1 0 10856 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_110
timestamp 1629484573
transform 1 0 11224 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_1  _518_
timestamp 1629484573
transform -1 0 12052 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_119
timestamp 1629484573
transform 1 0 12052 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _520_
timestamp 1629484573
transform 1 0 12788 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1629484573
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1629484573
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1629484573
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1629484573
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_147
timestamp 1629484573
transform 1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _413_
timestamp 1629484573
transform 1 0 14168 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _419_
timestamp 1629484573
transform 1 0 14996 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_159
timestamp 1629484573
transform 1 0 15732 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_163
timestamp 1629484573
transform 1 0 16100 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1629484573
transform -1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_11
timestamp 1629484573
transform 1 0 2116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1629484573
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1629484573
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _578_
timestamp 1629484573
transform 1 0 2208 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_19
timestamp 1629484573
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_34
timestamp 1629484573
transform 1 0 4232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1629484573
transform 1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1629484573
transform 1 0 4600 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 1629484573
transform 1 0 4876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _521_
timestamp 1629484573
transform 1 0 5244 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1629484573
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1629484573
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _488_
timestamp 1629484573
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_65
timestamp 1629484573
transform 1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_77
timestamp 1629484573
transform 1 0 8188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _540_
timestamp 1629484573
transform 1 0 7452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_84
timestamp 1629484573
transform 1 0 8832 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _403_
timestamp 1629484573
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _481_
timestamp 1629484573
transform -1 0 9476 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_91
timestamp 1629484573
transform 1 0 9476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1629484573
transform 1 0 10120 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _479_
timestamp 1629484573
transform -1 0 10948 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _480_
timestamp 1629484573
transform -1 0 10120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1629484573
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1629484573
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1629484573
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _477_
timestamp 1629484573
transform 1 0 11500 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_120
timestamp 1629484573
transform 1 0 12144 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _517_
timestamp 1629484573
transform 1 0 12512 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_9_129
timestamp 1629484573
transform 1 0 12972 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_135
timestamp 1629484573
transform 1 0 13524 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_139
timestamp 1629484573
transform 1 0 13892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _317_
timestamp 1629484573
transform -1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_145
timestamp 1629484573
transform 1 0 14444 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1629484573
transform 1 0 15180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _379_
timestamp 1629484573
transform -1 0 15180 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_160
timestamp 1629484573
transform 1 0 15824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1629484573
transform -1 0 16468 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1629484573
transform 1 0 15548 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1629484573
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1629484573
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1629484573
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _551_
timestamp 1629484573
transform 1 0 2484 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1629484573
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1629484573
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1629484573
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _550_
timestamp 1629484573
transform 1 0 4140 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_10_40
timestamp 1629484573
transform 1 0 4784 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_49
timestamp 1629484573
transform 1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1629484573
transform 1 0 5336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1629484573
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_63
timestamp 1629484573
transform 1 0 6900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _507_
timestamp 1629484573
transform 1 0 6624 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1629484573
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_72
timestamp 1629484573
transform 1 0 7728 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_76
timestamp 1629484573
transform 1 0 8096 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _506_
timestamp 1629484573
transform -1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _539_
timestamp 1629484573
transform -1 0 7728 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1629484573
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1629484573
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1629484573
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_1  _483_
timestamp 1629484573
transform 1 0 9292 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp 1629484573
transform 1 0 10028 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _505_
timestamp 1629484573
transform 1 0 10396 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_10_108
timestamp 1629484573
transform 1 0 11040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _482_
timestamp 1629484573
transform -1 0 11868 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_10_117
timestamp 1629484573
transform 1 0 11868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1629484573
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_128
timestamp 1629484573
transform 1 0 12880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1629484573
transform -1 0 12512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1629484573
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1629484573
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _356_
timestamp 1629484573
transform 1 0 14076 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _381_
timestamp 1629484573
transform 1 0 12972 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp 1629484573
transform 1 0 14720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _382_
timestamp 1629484573
transform 1 0 15088 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_10_157
timestamp 1629484573
transform 1 0 15548 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_163
timestamp 1629484573
transform 1 0 16100 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1629484573
transform -1 0 16468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1629484573
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1629484573
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1629484573
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _579_
timestamp 1629484573
transform -1 0 2116 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_11_23
timestamp 1629484573
transform 1 0 3220 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _552_
timestamp 1629484573
transform -1 0 3220 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_31
timestamp 1629484573
transform 1 0 3956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _522_
timestamp 1629484573
transform 1 0 4048 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_40
timestamp 1629484573
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _489_
timestamp 1629484573
transform 1 0 5152 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1629484573
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1629484573
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_61
timestamp 1629484573
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1629484573
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _357_
timestamp 1629484573
transform 1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_66
timestamp 1629484573
transform 1 0 7176 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 1629484573
transform 1 0 7912 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _508_
timestamp 1629484573
transform 1 0 8004 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_83
timestamp 1629484573
transform 1 0 8740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1629484573
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_92
timestamp 1629484573
transform 1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _478_
timestamp 1629484573
transform 1 0 9936 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1629484573
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1629484573
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1629484573
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1629484573
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  _355_
timestamp 1629484573
transform 1 0 11684 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_124
timestamp 1629484573
transform 1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _358_
timestamp 1629484573
transform 1 0 12880 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_11_135
timestamp 1629484573
transform 1 0 13524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _376_
timestamp 1629484573
transform 1 0 14076 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_11_146
timestamp 1629484573
transform 1 0 14536 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _383_
timestamp 1629484573
transform 1 0 14904 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_158
timestamp 1629484573
transform 1 0 15640 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1629484573
transform -1 0 16468 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_12
timestamp 1629484573
transform 1 0 2208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1629484573
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1629484573
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _580_
timestamp 1629484573
transform 1 0 1748 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1629484573
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output17
timestamp 1629484573
transform -1 0 2944 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1629484573
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_38
timestamp 1629484573
transform 1 0 4600 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1629484573
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _523_
timestamp 1629484573
transform 1 0 3864 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_50
timestamp 1629484573
transform 1 0 5704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_58
timestamp 1629484573
transform 1 0 6440 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_63
timestamp 1629484573
transform 1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _509_
timestamp 1629484573
transform -1 0 6900 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_75
timestamp 1629484573
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _511_
timestamp 1629484573
transform 1 0 7268 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1629484573
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1629484573
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _316_
timestamp 1629484573
transform 1 0 8924 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_12_101
timestamp 1629484573
transform 1 0 10396 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_95
timestamp 1629484573
transform 1 0 9844 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1629484573
transform 1 0 10488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_105
timestamp 1629484573
transform 1 0 10764 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _441_
timestamp 1629484573
transform 1 0 11132 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_12_116
timestamp 1629484573
transform 1 0 11776 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_124
timestamp 1629484573
transform 1 0 12512 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _322_
timestamp 1629484573
transform 1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_130
timestamp 1629484573
transform 1 0 13064 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1629484573
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1629484573
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _359_
timestamp 1629484573
transform 1 0 13156 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _375_
timestamp 1629484573
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_149
timestamp 1629484573
transform 1 0 14812 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_155
timestamp 1629484573
transform 1 0 15364 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_160
timestamp 1629484573
transform 1 0 15824 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1629484573
transform -1 0 16468 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1629484573
transform -1 0 15824 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1629484573
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1629484573
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_12
timestamp 1629484573
transform 1 0 2208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1629484573
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1629484573
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1629484573
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _581_
timestamp 1629484573
transform -1 0 2300 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _583_
timestamp 1629484573
transform -1 0 2208 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1629484573
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_21
timestamp 1629484573
transform 1 0 3036 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1629484573
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _555_
timestamp 1629484573
transform -1 0 3312 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _603_
timestamp 1629484573
transform -1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_33
timestamp 1629484573
transform 1 0 4140 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_34
timestamp 1629484573
transform 1 0 4232 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1629484573
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _554_
timestamp 1629484573
transform 1 0 3772 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_13_41
timestamp 1629484573
transform 1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 1629484573
transform 1 0 5336 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _456_
timestamp 1629484573
transform 1 0 5152 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _490_
timestamp 1629484573
transform 1 0 5428 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1629484573
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1629484573
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_54
timestamp 1629484573
transform 1 0 6072 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_62
timestamp 1629484573
transform 1 0 6808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1629484573
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _510_
timestamp 1629484573
transform 1 0 6900 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_13_73
timestamp 1629484573
transform 1 0 7820 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_68
timestamp 1629484573
transform 1 0 7360 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _473_
timestamp 1629484573
transform 1 0 7728 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _533_
timestamp 1629484573
transform 1 0 7084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_82
timestamp 1629484573
transform 1 0 8648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_89
timestamp 1629484573
transform 1 0 9292 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1629484573
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_88
timestamp 1629484573
transform 1 0 9200 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1629484573
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _333_
timestamp 1629484573
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _389_
timestamp 1629484573
transform 1 0 9016 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 1629484573
transform -1 0 8648 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_100
timestamp 1629484573
transform 1 0 10304 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_101
timestamp 1629484573
transform 1 0 10396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _410_
timestamp 1629484573
transform -1 0 10396 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _442_
timestamp 1629484573
transform -1 0 10304 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_13_104
timestamp 1629484573
transform 1 0 10672 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1629484573
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1629484573
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_110
timestamp 1629484573
transform 1 0 11224 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1629484573
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1629484573
transform 1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _346_
timestamp 1629484573
transform 1 0 11684 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _443_
timestamp 1629484573
transform 1 0 10764 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_13_124
timestamp 1629484573
transform 1 0 12512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_116
timestamp 1629484573
transform 1 0 11776 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_121
timestamp 1629484573
transform 1 0 12236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_125
timestamp 1629484573
transform 1 0 12604 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__and4_1  _334_
timestamp 1629484573
transform 1 0 12696 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _340_
timestamp 1629484573
transform 1 0 11868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _380_
timestamp 1629484573
transform -1 0 13156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_131
timestamp 1629484573
transform 1 0 13156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1629484573
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1629484573
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1629484573
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _353_
timestamp 1629484573
transform 1 0 14076 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _360_
timestamp 1629484573
transform 1 0 13524 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_143
timestamp 1629484573
transform 1 0 14260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_146
timestamp 1629484573
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_150
timestamp 1629484573
transform 1 0 14904 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  _320_
timestamp 1629484573
transform 1 0 14996 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _420_
timestamp 1629484573
transform 1 0 14628 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_155
timestamp 1629484573
transform 1 0 15364 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_163
timestamp 1629484573
transform 1 0 16100 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_160
timestamp 1629484573
transform 1 0 15824 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1629484573
transform -1 0 16468 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1629484573
transform -1 0 16468 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1629484573
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1629484573
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _582_
timestamp 1629484573
transform -1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1629484573
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_20
timestamp 1629484573
transform 1 0 2944 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _602_
timestamp 1629484573
transform 1 0 2668 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_28
timestamp 1629484573
transform 1 0 3680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_37
timestamp 1629484573
transform 1 0 4508 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _524_
timestamp 1629484573
transform 1 0 3864 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1629484573
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _491_
timestamp 1629484573
transform 1 0 4876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1629484573
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1629484573
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_61
timestamp 1629484573
transform 1 0 6716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1629484573
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _474_
timestamp 1629484573
transform -1 0 6716 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_68
timestamp 1629484573
transform 1 0 7360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _471_
timestamp 1629484573
transform -1 0 7360 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _503_
timestamp 1629484573
transform 1 0 7728 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_15_82
timestamp 1629484573
transform 1 0 8648 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_88
timestamp 1629484573
transform 1 0 9200 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_1  _446_
timestamp 1629484573
transform 1 0 9292 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_97
timestamp 1629484573
transform 1 0 10028 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _390_
timestamp 1629484573
transform 1 0 10396 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1629484573
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1629484573
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _445_
timestamp 1629484573
transform -1 0 11960 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_15_118
timestamp 1629484573
transform 1 0 11960 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _318_
timestamp 1629484573
transform 1 0 12696 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_15_133
timestamp 1629484573
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_140
timestamp 1629484573
transform 1 0 13984 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _348_
timestamp 1629484573
transform -1 0 13984 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_148
timestamp 1629484573
transform 1 0 14720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_1  _632_
timestamp 1629484573
transform -1 0 15548 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_15_157
timestamp 1629484573
transform 1 0 15548 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_163
timestamp 1629484573
transform 1 0 16100 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1629484573
transform -1 0 16468 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1629484573
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1629484573
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _605_
timestamp 1629484573
transform 1 0 1656 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_13
timestamp 1629484573
transform 1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1629484573
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _553_
timestamp 1629484573
transform 1 0 2668 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1629484573
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_38
timestamp 1629484573
transform 1 0 4600 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1629484573
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _525_
timestamp 1629484573
transform 1 0 3864 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_50
timestamp 1629484573
transform 1 0 5704 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_59
timestamp 1629484573
transform 1 0 6532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _472_
timestamp 1629484573
transform -1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _476_
timestamp 1629484573
transform 1 0 6900 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_71
timestamp 1629484573
transform 1 0 7636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _475_
timestamp 1629484573
transform 1 0 8004 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1629484573
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1629484573
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp 1629484573
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1629484573
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_97
timestamp 1629484573
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _388_
timestamp 1629484573
transform -1 0 10672 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _470_
timestamp 1629484573
transform 1 0 9384 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_16_104
timestamp 1629484573
transform 1 0 10672 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_112
timestamp 1629484573
transform 1 0 11408 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _409_
timestamp 1629484573
transform 1 0 11500 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_120
timestamp 1629484573
transform 1 0 12144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_127
timestamp 1629484573
transform 1 0 12788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1629484573
transform -1 0 12788 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_134
timestamp 1629484573
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1629484573
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _326_
timestamp 1629484573
transform 1 0 13156 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _335_
timestamp 1629484573
transform 1 0 14076 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1629484573
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_160
timestamp 1629484573
transform 1 0 15824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1629484573
transform -1 0 16468 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  _633_
timestamp 1629484573
transform -1 0 15824 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1629484573
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1629484573
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1629484573
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _604_
timestamp 1629484573
transform 1 0 1840 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1629484573
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _526_
timestamp 1629484573
transform 1 0 2852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1629484573
transform 1 0 3588 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _492_
timestamp 1629484573
transform 1 0 3956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_39
timestamp 1629484573
transform 1 0 4692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 1629484573
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _457_
timestamp 1629484573
transform 1 0 5152 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1629484573
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1629484573
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1629484573
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _504_
timestamp 1629484573
transform 1 0 6900 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_71
timestamp 1629484573
transform 1 0 7636 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _438_
timestamp 1629484573
transform -1 0 8464 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_17_80
timestamp 1629484573
transform 1 0 8464 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1629484573
transform 1 0 9200 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _411_
timestamp 1629484573
transform 1 0 9292 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_17_94
timestamp 1629484573
transform 1 0 9752 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _385_
timestamp 1629484573
transform -1 0 11040 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1629484573
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1629484573
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1629484573
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _387_
timestamp 1629484573
transform -1 0 12236 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_17_121
timestamp 1629484573
transform 1 0 12236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_128
timestamp 1629484573
transform 1 0 12880 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1629484573
transform -1 0 12880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_136
timestamp 1629484573
transform 1 0 13616 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _327_
timestamp 1629484573
transform -1 0 14352 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_17_144
timestamp 1629484573
transform 1 0 14352 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_152
timestamp 1629484573
transform 1 0 15088 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _367_
timestamp 1629484573
transform 1 0 15180 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1629484573
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_163
timestamp 1629484573
transform 1 0 16100 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1629484573
transform -1 0 16468 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1629484573
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1629484573
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _558_
timestamp 1629484573
transform 1 0 1564 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_13
timestamp 1629484573
transform 1 0 2300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1629484573
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _556_
timestamp 1629484573
transform -1 0 2944 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1629484573
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1629484573
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1629484573
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1629484573
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_65
timestamp 1629484573
transform 1 0 7084 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_73
timestamp 1629484573
transform 1 0 7820 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _402_
timestamp 1629484573
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _468_
timestamp 1629484573
transform 1 0 7176 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1629484573
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1629484573
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1629484573
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o21ba_1  _437_
timestamp 1629484573
transform 1 0 9200 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_96
timestamp 1629484573
transform 1 0 9936 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _394_
timestamp 1629484573
transform -1 0 11224 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_18_110
timestamp 1629484573
transform 1 0 11224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _313_
timestamp 1629484573
transform -1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_117
timestamp 1629484573
transform 1 0 11868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_127
timestamp 1629484573
transform 1 0 12788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _350_
timestamp 1629484573
transform -1 0 12788 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1629484573
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1629484573
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _332_
timestamp 1629484573
transform 1 0 13156 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _336_
timestamp 1629484573
transform -1 0 14720 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1629484573
transform 1 0 14720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _366_
timestamp 1629484573
transform -1 0 15824 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_160
timestamp 1629484573
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1629484573
transform -1 0 16468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_11
timestamp 1629484573
transform 1 0 2116 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1629484573
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1629484573
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1629484573
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1629484573
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _528_
timestamp 1629484573
transform 1 0 2116 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output30
timestamp 1629484573
transform -1 0 2116 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_18
timestamp 1629484573
transform 1 0 2760 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_24
timestamp 1629484573
transform 1 0 3312 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_17
timestamp 1629484573
transform 1 0 2668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1629484573
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _495_
timestamp 1629484573
transform 1 0 3404 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _527_
timestamp 1629484573
transform 1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _557_
timestamp 1629484573
transform 1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_33
timestamp 1629484573
transform 1 0 4140 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_37
timestamp 1629484573
transform 1 0 4508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1629484573
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _494_
timestamp 1629484573
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_41
timestamp 1629484573
transform 1 0 4876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_41
timestamp 1629484573
transform 1 0 4876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_50
timestamp 1629484573
transform 1 0 5704 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_1  _459_
timestamp 1629484573
transform 1 0 5152 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _460_
timestamp 1629484573
transform 1 0 4968 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1629484573
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1629484573
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_62
timestamp 1629484573
transform 1 0 6808 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1629484573
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _440_
timestamp 1629484573
transform 1 0 6532 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_67
timestamp 1629484573
transform 1 0 7268 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_68
timestamp 1629484573
transform 1 0 7360 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_74
timestamp 1629484573
transform 1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _436_
timestamp 1629484573
transform -1 0 7912 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _439_
timestamp 1629484573
transform 1 0 7636 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_79
timestamp 1629484573
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_86
timestamp 1629484573
transform 1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1629484573
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1629484573
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _341_
timestamp 1629484573
transform 1 0 8740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _458_
timestamp 1629484573
transform 1 0 8924 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1629484573
transform 1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_92
timestamp 1629484573
transform 1 0 9568 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1629484573
transform 1 0 10304 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _408_
timestamp 1629484573
transform -1 0 10948 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _412_
timestamp 1629484573
transform 1 0 9384 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1629484573
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1629484573
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_103
timestamp 1629484573
transform 1 0 10580 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_114
timestamp 1629484573
transform 1 0 11592 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1629484573
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _395_
timestamp 1629484573
transform 1 0 11500 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _400_
timestamp 1629484573
transform 1 0 10948 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_19_118
timestamp 1629484573
transform 1 0 11960 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_124
timestamp 1629484573
transform 1 0 12512 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_123
timestamp 1629484573
transform 1 0 12420 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _349_
timestamp 1629484573
transform -1 0 13248 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _391_
timestamp 1629484573
transform 1 0 11960 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_19_132
timestamp 1629484573
transform 1 0 13248 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1629484573
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1629484573
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _314_
timestamp 1629484573
transform 1 0 13984 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _328_
timestamp 1629484573
transform 1 0 14076 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _342_
timestamp 1629484573
transform 1 0 13156 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_19_145
timestamp 1629484573
transform 1 0 14444 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_146
timestamp 1629484573
transform 1 0 14536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _337_
timestamp 1629484573
transform 1 0 14904 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _338_
timestamp 1629484573
transform 1 0 14996 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_159
timestamp 1629484573
transform 1 0 15732 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_163
timestamp 1629484573
transform 1 0 16100 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_155
timestamp 1629484573
transform 1 0 15364 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_163
timestamp 1629484573
transform 1 0 16100 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1629484573
transform -1 0 16468 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1629484573
transform -1 0 16468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_6
timestamp 1629484573
transform 1 0 1656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1629484573
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1629484573
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _532_
timestamp 1629484573
transform 1 0 2024 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_18
timestamp 1629484573
transform 1 0 2760 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _502_
timestamp 1629484573
transform 1 0 3312 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_21_31
timestamp 1629484573
transform 1 0 3956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_39
timestamp 1629484573
transform 1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_48
timestamp 1629484573
transform 1 0 5520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _493_
timestamp 1629484573
transform 1 0 4876 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_21_57
timestamp 1629484573
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1629484573
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_65
timestamp 1629484573
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_70
timestamp 1629484573
transform 1 0 7544 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_77
timestamp 1629484573
transform 1 0 8188 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _405_
timestamp 1629484573
transform 1 0 7912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _407_
timestamp 1629484573
transform -1 0 7544 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _421_
timestamp 1629484573
transform 1 0 9292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_97
timestamp 1629484573
transform 1 0 10028 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1629484573
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1629484573
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1629484573
transform -1 0 11040 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _396_
timestamp 1629484573
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_121
timestamp 1629484573
transform 1 0 12236 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_128
timestamp 1629484573
transform 1 0 12880 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1629484573
transform -1 0 12880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_136
timestamp 1629484573
transform 1 0 13616 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o21ba_1  _352_
timestamp 1629484573
transform 1 0 13708 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_145
timestamp 1629484573
transform 1 0 14444 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_153
timestamp 1629484573
transform 1 0 15180 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_1  _634_
timestamp 1629484573
transform 1 0 15272 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_160
timestamp 1629484573
transform 1 0 15824 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1629484573
transform -1 0 16468 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_10
timestamp 1629484573
transform 1 0 2024 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1629484573
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1629484573
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1629484573
transform 1 0 1748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1629484573
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _499_
timestamp 1629484573
transform 1 0 2760 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1629484573
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp 1629484573
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1629484573
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _496_
timestamp 1629484573
transform 1 0 4232 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1629484573
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1629484573
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_72
timestamp 1629484573
transform 1 0 7728 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _406_
timestamp 1629484573
transform 1 0 8096 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _461_
timestamp 1629484573
transform 1 0 7084 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1629484573
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1629484573
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1629484573
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _422_
timestamp 1629484573
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_101
timestamp 1629484573
transform 1 0 10396 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_93
timestamp 1629484573
transform 1 0 9660 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_107
timestamp 1629484573
transform 1 0 10948 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _423_
timestamp 1629484573
transform 1 0 11316 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _631_
timestamp 1629484573
transform 1 0 10672 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_118
timestamp 1629484573
transform 1 0 11960 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _384_
timestamp 1629484573
transform 1 0 12328 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_130
timestamp 1629484573
transform 1 0 13064 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1629484573
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp 1629484573
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1629484573
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_150
timestamp 1629484573
transform 1 0 14904 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_154
timestamp 1629484573
transform 1 0 15272 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _329_
timestamp 1629484573
transform -1 0 14904 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_160
timestamp 1629484573
transform 1 0 15824 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1629484573
transform -1 0 16468 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _368_
timestamp 1629484573
transform -1 0 15824 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1629484573
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp 1629484573
transform 1 0 1932 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1629484573
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _530_
timestamp 1629484573
transform -1 0 2760 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_18
timestamp 1629484573
transform 1 0 2760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_25
timestamp 1629484573
transform 1 0 3404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _498_
timestamp 1629484573
transform -1 0 3404 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_37
timestamp 1629484573
transform 1 0 4508 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _463_
timestamp 1629484573
transform 1 0 3772 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_49
timestamp 1629484573
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _462_
timestamp 1629484573
transform 1 0 4876 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1629484573
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 1629484573
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1629484573
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _425_
timestamp 1629484573
transform 1 0 6440 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_66
timestamp 1629484573
transform 1 0 7176 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_72
timestamp 1629484573
transform 1 0 7728 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _424_
timestamp 1629484573
transform 1 0 7820 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1629484573
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1629484573
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1629484573
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1629484573
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1629484573
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _397_
timestamp 1629484573
transform -1 0 12236 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_121
timestamp 1629484573
transform 1 0 12236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_128
timestamp 1629484573
transform 1 0 12880 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _331_
timestamp 1629484573
transform 1 0 12604 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _344_
timestamp 1629484573
transform 1 0 13616 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_143
timestamp 1629484573
transform 1 0 14260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _343_
timestamp 1629484573
transform -1 0 15364 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_155
timestamp 1629484573
transform 1 0 15364 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_163
timestamp 1629484573
transform 1 0 16100 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1629484573
transform -1 0 16468 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1629484573
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_8
timestamp 1629484573
transform 1 0 1840 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1629484573
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _531_
timestamp 1629484573
transform -1 0 1840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_18
timestamp 1629484573
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _529_
timestamp 1629484573
transform 1 0 2392 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1629484573
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_34
timestamp 1629484573
transform 1 0 4232 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1629484573
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _497_
timestamp 1629484573
transform -1 0 4232 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_24_46
timestamp 1629484573
transform 1 0 5336 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_58
timestamp 1629484573
transform 1 0 6440 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_70
timestamp 1629484573
transform 1 0 7544 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1629484573
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1629484573
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1629484573
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1629484573
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_98
timestamp 1629484573
transform 1 0 10120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _363_
timestamp 1629484573
transform -1 0 10948 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1629484573
transform 1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_107
timestamp 1629484573
transform 1 0 10948 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_111
timestamp 1629484573
transform 1 0 11316 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1629484573
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1629484573
transform -1 0 11684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_122
timestamp 1629484573
transform 1 0 12328 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _351_
timestamp 1629484573
transform 1 0 12696 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1629484573
transform 1 0 12052 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_132
timestamp 1629484573
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1629484573
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1629484573
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1629484573
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_154
timestamp 1629484573
transform 1 0 15272 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _369_
timestamp 1629484573
transform -1 0 15272 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_162
timestamp 1629484573
transform 1 0 16008 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1629484573
transform -1 0 16468 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1629484573
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1629484573
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_15
timestamp 1629484573
transform 1 0 2484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_23
timestamp 1629484573
transform 1 0 3220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_33
timestamp 1629484573
transform 1 0 4140 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _500_
timestamp 1629484573
transform 1 0 3496 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_25_39
timestamp 1629484573
transform 1 0 4692 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_43
timestamp 1629484573
transform 1 0 5060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _426_
timestamp 1629484573
transform -1 0 5888 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _464_
timestamp 1629484573
transform 1 0 4784 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1629484573
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1629484573
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1629484573
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _466_
timestamp 1629484573
transform 1 0 6532 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_25_66
timestamp 1629484573
transform 1 0 7176 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2oi_1  _433_
timestamp 1629484573
transform 1 0 7728 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_25_79
timestamp 1629484573
transform 1 0 8372 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_87
timestamp 1629484573
transform 1 0 9108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _371_
timestamp 1629484573
transform -1 0 9660 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1629484573
transform 1 0 9660 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_97
timestamp 1629484573
transform 1 0 10028 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_1  _365_
timestamp 1629484573
transform 1 0 10120 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_104
timestamp 1629484573
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1629484573
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _429_
timestamp 1629484573
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_121
timestamp 1629484573
transform 1 0 12236 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_137
timestamp 1629484573
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _362_
timestamp 1629484573
transform 1 0 12972 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_149
timestamp 1629484573
transform 1 0 14812 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _635_
timestamp 1629484573
transform -1 0 15732 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output25
timestamp 1629484573
transform 1 0 14444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1629484573
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_163
timestamp 1629484573
transform 1 0 16100 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1629484573
transform -1 0 16468 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1629484573
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_9
timestamp 1629484573
transform 1 0 1932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_11
timestamp 1629484573
transform 1 0 2116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1629484573
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1629484573
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1629484573
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _501_
timestamp 1629484573
transform 1 0 2024 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1629484573
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_17
timestamp 1629484573
transform 1 0 2668 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp 1629484573
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_19
timestamp 1629484573
transform 1 0 2852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output18
timestamp 1629484573
transform -1 0 2852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_36
timestamp 1629484573
transform 1 0 4416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1629484573
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_29
timestamp 1629484573
transform 1 0 3772 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_37
timestamp 1629484573
transform 1 0 4508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1629484573
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1629484573
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _467_
timestamp 1629484573
transform -1 0 4416 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output22
timestamp 1629484573
transform -1 0 4508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1629484573
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1629484573
transform 1 0 5244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1629484573
transform 1 0 5612 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _428_
timestamp 1629484573
transform -1 0 6348 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _465_
timestamp 1629484573
transform -1 0 5428 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output31
timestamp 1629484573
transform -1 0 5244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_57
timestamp 1629484573
transform 1 0 6348 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1629484573
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1629484573
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _431_
timestamp 1629484573
transform -1 0 7636 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1629484573
transform 1 0 6348 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_26_71
timestamp 1629484573
transform 1 0 7636 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_75
timestamp 1629484573
transform 1 0 8004 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_67
timestamp 1629484573
transform 1 0 7268 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _373_
timestamp 1629484573
transform 1 0 8096 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output27
timestamp 1629484573
transform -1 0 8372 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1629484573
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1629484573
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_79
timestamp 1629484573
transform 1 0 8372 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_83
timestamp 1629484573
transform 1 0 8740 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_85
timestamp 1629484573
transform 1 0 8924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1629484573
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1629484573
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _430_
timestamp 1629484573
transform -1 0 9476 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _432_
timestamp 1629484573
transform -1 0 9476 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_26_91
timestamp 1629484573
transform 1 0 9476 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_101
timestamp 1629484573
transform 1 0 10396 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_91
timestamp 1629484573
transform 1 0 9476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_95
timestamp 1629484573
transform 1 0 9844 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _629_
timestamp 1629484573
transform 1 0 9936 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _630_
timestamp 1629484573
transform -1 0 10580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_103
timestamp 1629484573
transform 1 0 10580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_111
timestamp 1629484573
transform 1 0 11316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1629484573
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1629484573
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1629484573
transform 1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _398_
timestamp 1629484573
transform -1 0 12236 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _399_
timestamp 1629484573
transform 1 0 11500 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_26_121
timestamp 1629484573
transform 1 0 12236 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_127
timestamp 1629484573
transform 1 0 12788 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_120
timestamp 1629484573
transform 1 0 12144 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_128
timestamp 1629484573
transform 1 0 12880 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _361_
timestamp 1629484573
transform 1 0 12880 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output28
timestamp 1629484573
transform -1 0 12880 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1629484573
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_135
timestamp 1629484573
transform 1 0 13524 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_139
timestamp 1629484573
transform 1 0 13892 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1629484573
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1629484573
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _374_
timestamp 1629484573
transform -1 0 14720 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1629484573
transform -1 0 14352 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1629484573
transform -1 0 13524 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1629484573
transform 1 0 14720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1629484573
transform 1 0 15088 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_144
timestamp 1629484573
transform 1 0 14352 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_148
timestamp 1629484573
transform 1 0 14720 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_152
timestamp 1629484573
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _370_
timestamp 1629484573
transform 1 0 15180 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1629484573
transform -1 0 15088 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_158
timestamp 1629484573
transform 1 0 15640 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_160
timestamp 1629484573
transform 1 0 15824 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1629484573
transform -1 0 16468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1629484573
transform -1 0 16468 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output26
timestamp 1629484573
transform 1 0 15456 0 -1 17408
box -38 -48 406 592
<< labels >>
rlabel metal2 s 17498 18928 17554 19728 4 A[0]
port 1 nsew
rlabel metal3 s 0 17144 800 17264 4 A[1]
port 2 nsew
rlabel metal3 s 0 5720 800 5840 4 A[2]
port 3 nsew
rlabel metal2 s 7746 0 7802 800 4 A[3]
port 4 nsew
rlabel metal2 s 5906 18928 5962 19728 4 A[4]
port 5 nsew
rlabel metal2 s 11794 18928 11850 19728 4 A[5]
port 6 nsew
rlabel metal2 s 13450 0 13506 800 4 A[6]
port 7 nsew
rlabel metal3 s 16784 8168 17584 8288 4 A[7]
port 8 nsew
rlabel metal2 s 11610 0 11666 800 4 B[0]
port 9 nsew
rlabel metal3 s 16784 11160 17584 11280 4 B[1]
port 10 nsew
rlabel metal3 s 0 2728 800 2848 4 B[2]
port 11 nsew
rlabel metal2 s 18 0 74 800 4 B[3]
port 12 nsew
rlabel metal2 s 13634 18928 13690 19728 4 B[4]
port 13 nsew
rlabel metal2 s 15658 18928 15714 19728 4 B[5]
port 14 nsew
rlabel metal3 s 0 14152 800 14272 4 B[6]
port 15 nsew
rlabel metal2 s 17498 0 17554 800 4 B[7]
port 16 nsew
rlabel metal3 s 0 8440 800 8560 4 M[0]
port 17 nsew
rlabel metal2 s 18 18928 74 19728 4 M[10]
port 18 nsew
rlabel metal2 s 15474 0 15530 800 4 M[11]
port 19 nsew
rlabel metal2 s 1858 0 1914 800 4 M[12]
port 20 nsew
rlabel metal2 s 3882 0 3938 800 4 M[13]
port 21 nsew
rlabel metal2 s 4066 18928 4122 19728 4 M[14]
port 22 nsew
rlabel metal3 s 16784 2456 17584 2576 4 M[15]
port 23 nsew
rlabel metal2 s 5722 0 5778 800 4 M[1]
port 24 nsew
rlabel metal3 s 16784 13880 17584 14000 4 M[2]
port 25 nsew
rlabel metal3 s 16784 16872 17584 16992 4 M[3]
port 26 nsew
rlabel metal2 s 7930 18928 7986 19728 4 M[4]
port 27 nsew
rlabel metal2 s 9770 18928 9826 19728 4 M[5]
port 28 nsew
rlabel metal2 s 9586 0 9642 800 4 M[6]
port 29 nsew
rlabel metal3 s 0 11432 800 11552 4 M[7]
port 30 nsew
rlabel metal2 s 2042 18928 2098 19728 4 M[8]
port 31 nsew
rlabel metal3 s 16784 5448 17584 5568 4 M[9]
port 32 nsew
rlabel metal5 s 1104 7046 16468 7366 4 VGND
port 33 nsew
rlabel metal5 s 1104 4506 16468 4826 4 VPWR
port 34 nsew
<< properties >>
string FIXED_BBOX 0 0 17584 19728
<< end >>
